module fpgasoc_fetal_ecg();


endmodule
