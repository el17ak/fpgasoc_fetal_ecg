// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition"

// DATE "05/10/2022 21:57:12"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Computer_System (
	hps_f2h_irq0_irq,
	hps_io_hps_io_emac1_inst_TX_CLK,
	hps_io_hps_io_emac1_inst_TXD0,
	hps_io_hps_io_emac1_inst_TXD1,
	hps_io_hps_io_emac1_inst_TXD2,
	hps_io_hps_io_emac1_inst_TXD3,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_MDIO,
	hps_io_hps_io_emac1_inst_MDC,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_emac1_inst_TX_CTL,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_qspi_inst_IO0,
	hps_io_hps_io_qspi_inst_IO1,
	hps_io_hps_io_qspi_inst_IO2,
	hps_io_hps_io_qspi_inst_IO3,
	hps_io_hps_io_qspi_inst_SS0,
	hps_io_hps_io_qspi_inst_CLK,
	hps_io_hps_io_sdio_inst_CMD,
	hps_io_hps_io_sdio_inst_D0,
	hps_io_hps_io_sdio_inst_D1,
	hps_io_hps_io_sdio_inst_CLK,
	hps_io_hps_io_sdio_inst_D2,
	hps_io_hps_io_sdio_inst_D3,
	hps_io_hps_io_usb1_inst_D0,
	hps_io_hps_io_usb1_inst_D1,
	hps_io_hps_io_usb1_inst_D2,
	hps_io_hps_io_usb1_inst_D3,
	hps_io_hps_io_usb1_inst_D4,
	hps_io_hps_io_usb1_inst_D5,
	hps_io_hps_io_usb1_inst_D6,
	hps_io_hps_io_usb1_inst_D7,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_STP,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	hps_io_hps_io_spim1_inst_CLK,
	hps_io_hps_io_spim1_inst_MOSI,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_spim1_inst_SS0,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_uart0_inst_TX,
	hps_io_hps_io_i2c0_inst_SDA,
	hps_io_hps_io_i2c0_inst_SCL,
	hps_io_hps_io_i2c1_inst_SDA,
	hps_io_hps_io_i2c1_inst_SCL,
	hps_io_hps_io_gpio_inst_GPIO09,
	hps_io_hps_io_gpio_inst_GPIO35,
	hps_io_hps_io_gpio_inst_GPIO40,
	hps_io_hps_io_gpio_inst_GPIO41,
	hps_io_hps_io_gpio_inst_GPIO48,
	hps_io_hps_io_gpio_inst_GPIO53,
	hps_io_hps_io_gpio_inst_GPIO54,
	hps_io_hps_io_gpio_inst_GPIO61,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	onchip_sram_clk2_clk,
	onchip_sram_reset2_reset,
	onchip_sram_reset2_reset_req,
	onchip_sram_s2_address,
	onchip_sram_s2_chipselect,
	onchip_sram_s2_clken,
	onchip_sram_s2_write,
	onchip_sram_s2_readdata,
	onchip_sram_s2_writedata,
	onchip_sram_s2_byteenable,
	sdram_clk_clk,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset)/* synthesis synthesis_greybox=0 */;
input 	[31:0] hps_f2h_irq0_irq;
output 	hps_io_hps_io_emac1_inst_TX_CLK;
output 	hps_io_hps_io_emac1_inst_TXD0;
output 	hps_io_hps_io_emac1_inst_TXD1;
output 	hps_io_hps_io_emac1_inst_TXD2;
output 	hps_io_hps_io_emac1_inst_TXD3;
input 	hps_io_hps_io_emac1_inst_RXD0;
inout 	hps_io_hps_io_emac1_inst_MDIO;
output 	hps_io_hps_io_emac1_inst_MDC;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
output 	hps_io_hps_io_emac1_inst_TX_CTL;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
inout 	hps_io_hps_io_qspi_inst_IO0;
inout 	hps_io_hps_io_qspi_inst_IO1;
inout 	hps_io_hps_io_qspi_inst_IO2;
inout 	hps_io_hps_io_qspi_inst_IO3;
output 	hps_io_hps_io_qspi_inst_SS0;
output 	hps_io_hps_io_qspi_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_CMD;
inout 	hps_io_hps_io_sdio_inst_D0;
inout 	hps_io_hps_io_sdio_inst_D1;
output 	hps_io_hps_io_sdio_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_D2;
inout 	hps_io_hps_io_sdio_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D0;
inout 	hps_io_hps_io_usb1_inst_D1;
inout 	hps_io_hps_io_usb1_inst_D2;
inout 	hps_io_hps_io_usb1_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D4;
inout 	hps_io_hps_io_usb1_inst_D5;
inout 	hps_io_hps_io_usb1_inst_D6;
inout 	hps_io_hps_io_usb1_inst_D7;
input 	hps_io_hps_io_usb1_inst_CLK;
output 	hps_io_hps_io_usb1_inst_STP;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
output 	hps_io_hps_io_spim1_inst_CLK;
output 	hps_io_hps_io_spim1_inst_MOSI;
input 	hps_io_hps_io_spim1_inst_MISO;
output 	hps_io_hps_io_spim1_inst_SS0;
input 	hps_io_hps_io_uart0_inst_RX;
output 	hps_io_hps_io_uart0_inst_TX;
inout 	hps_io_hps_io_i2c0_inst_SDA;
inout 	hps_io_hps_io_i2c0_inst_SCL;
inout 	hps_io_hps_io_i2c1_inst_SDA;
inout 	hps_io_hps_io_i2c1_inst_SCL;
inout 	hps_io_hps_io_gpio_inst_GPIO09;
inout 	hps_io_hps_io_gpio_inst_GPIO35;
inout 	hps_io_hps_io_gpio_inst_GPIO40;
inout 	hps_io_hps_io_gpio_inst_GPIO41;
inout 	hps_io_hps_io_gpio_inst_GPIO48;
inout 	hps_io_hps_io_gpio_inst_GPIO53;
inout 	hps_io_hps_io_gpio_inst_GPIO54;
inout 	hps_io_hps_io_gpio_inst_GPIO61;
output 	[14:0] memory_mem_a;
output 	[2:0] memory_mem_ba;
output 	memory_mem_ck;
output 	memory_mem_ck_n;
output 	memory_mem_cke;
output 	memory_mem_cs_n;
output 	memory_mem_ras_n;
output 	memory_mem_cas_n;
output 	memory_mem_we_n;
output 	memory_mem_reset_n;
inout 	[31:0] memory_mem_dq;
inout 	[3:0] memory_mem_dqs;
inout 	[3:0] memory_mem_dqs_n;
output 	memory_mem_odt;
output 	[3:0] memory_mem_dm;
input 	memory_oct_rzqin;
input 	onchip_sram_clk2_clk;
input 	onchip_sram_reset2_reset;
input 	onchip_sram_reset2_reset_req;
input 	[13:0] onchip_sram_s2_address;
input 	onchip_sram_s2_chipselect;
input 	onchip_sram_s2_clken;
input 	onchip_sram_s2_write;
output 	[31:0] onchip_sram_s2_readdata;
input 	[31:0] onchip_sram_s2_writedata;
input 	[3:0] onchip_sram_s2_byteenable;
output 	sdram_clk_clk;
input 	system_pll_ref_clk_clk;
input 	system_pll_ref_reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_ARREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_AWREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_BVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_WREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[0] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[1] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[2] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[3] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[4] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[5] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[6] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[7] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[8] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[9] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[10] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[11] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[12] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[13] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[14] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[15] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[16] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[17] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[18] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[19] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[20] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[21] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[22] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[23] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[24] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[25] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[26] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[27] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[28] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[29] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[30] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[31] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[32] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[33] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[34] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[35] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[36] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[37] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[38] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[39] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[40] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[41] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[42] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[43] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[44] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[45] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[46] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[47] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[48] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[49] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[50] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[51] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[52] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[53] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[54] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[55] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[56] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[57] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[58] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[59] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[60] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[61] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[62] ;
wire \arm_a9_hps|fpga_interfaces|f2h_RDATA[63] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_BREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_RREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WLAST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[12] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[13] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[14] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[15] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[16] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[17] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[18] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[19] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[20] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[21] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[22] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[23] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[24] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[25] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[26] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[27] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[28] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[29] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[30] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[31] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[3] ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a32~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a0~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a33~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a1~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a34~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a2~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a35~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a3~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a36~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a4~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a37~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a5~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a38~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a6~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a39~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a7~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a40~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a8~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a41~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a9~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a42~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a10~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a43~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a11~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a44~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a12~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a45~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a13~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a46~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a14~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a47~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a15~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a56~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a24~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a57~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a25~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a58~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a26~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a59~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a27~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a60~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a28~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a61~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a29~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a62~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a30~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a63~portadataout ;
wire \onchip_sram|the_altsyncram|auto_generated|ram_block1a31~portadataout ;
wire \system_pll|sys_pll|altera_pll_i|outclk_wire[1] ;
wire \system_pll|sys_pll|altera_pll_i|outclk_wire[0] ;
wire \system_pll|sys_pll|altera_pll_i|locked_wire[0] ;
wire \dma_1|readaddress[2]~q ;
wire \dma_1|readaddress[3]~q ;
wire \dma_1|readaddress[4]~q ;
wire \dma_1|readaddress[5]~q ;
wire \dma_1|readaddress[6]~q ;
wire \dma_1|readaddress[7]~q ;
wire \dma_1|readaddress[8]~q ;
wire \dma_1|readaddress[9]~q ;
wire \dma_1|readaddress[10]~q ;
wire \dma_1|readaddress[11]~q ;
wire \dma_1|readaddress[12]~q ;
wire \dma_1|readaddress[13]~q ;
wire \dma_1|readaddress[14]~q ;
wire \dma_1|readaddress[15]~q ;
wire \dma_1|readaddress[16]~q ;
wire \dma_1|readaddress[17]~q ;
wire \dma_1|readaddress[18]~q ;
wire \dma_1|readaddress[19]~q ;
wire \dma_1|readaddress[20]~q ;
wire \dma_1|readaddress[21]~q ;
wire \dma_1|readaddress[22]~q ;
wire \dma_1|readaddress[23]~q ;
wire \dma_1|readaddress[24]~q ;
wire \dma_1|readaddress[25]~q ;
wire \dma_1|readaddress[26]~q ;
wire \dma_1|readaddress[27]~q ;
wire \dma_1|readaddress[28]~q ;
wire \dma_1|readaddress[29]~q ;
wire \dma_1|readaddress[30]~q ;
wire \dma_1|readaddress[31]~q ;
wire \dma_2|writeaddress[2]~q ;
wire \dma_2|writeaddress[3]~q ;
wire \dma_2|writeaddress[4]~q ;
wire \dma_2|writeaddress[5]~q ;
wire \dma_2|writeaddress[6]~q ;
wire \dma_2|writeaddress[7]~q ;
wire \dma_2|writeaddress[8]~q ;
wire \dma_2|writeaddress[9]~q ;
wire \dma_2|writeaddress[10]~q ;
wire \dma_2|writeaddress[11]~q ;
wire \dma_2|writeaddress[12]~q ;
wire \dma_2|writeaddress[13]~q ;
wire \dma_2|writeaddress[14]~q ;
wire \dma_2|writeaddress[15]~q ;
wire \dma_2|writeaddress[16]~q ;
wire \dma_2|writeaddress[17]~q ;
wire \dma_2|writeaddress[18]~q ;
wire \dma_2|writeaddress[19]~q ;
wire \dma_2|writeaddress[20]~q ;
wire \dma_2|writeaddress[21]~q ;
wire \dma_2|writeaddress[22]~q ;
wire \dma_2|writeaddress[23]~q ;
wire \dma_2|writeaddress[24]~q ;
wire \dma_2|writeaddress[25]~q ;
wire \dma_2|writeaddress[26]~q ;
wire \dma_2|writeaddress[27]~q ;
wire \dma_2|writeaddress[28]~q ;
wire \dma_2|writeaddress[29]~q ;
wire \dma_2|writeaddress[30]~q ;
wire \dma_2|writeaddress[31]~q ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[0] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[1] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[2] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[3] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[4] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[5] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[6] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[7] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[8] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[9] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[10] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[11] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[12] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[13] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[14] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[15] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[16] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[17] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[18] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[19] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[20] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[21] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[22] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[23] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[24] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[25] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[26] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[27] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[28] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[29] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[30] ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[31] ;
wire \dma_2|writeaddress[1]~q ;
wire \dma_2|writeaddress[0]~q ;
wire \dma_2|readaddress[15]~q ;
wire \dma_1|writeaddress[15]~q ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[0] ;
wire \dma_2|readaddress[2]~q ;
wire \dma_1|writeaddress[2]~q ;
wire \dma_2|readaddress[3]~q ;
wire \dma_1|writeaddress[3]~q ;
wire \dma_2|readaddress[4]~q ;
wire \dma_1|writeaddress[4]~q ;
wire \dma_2|readaddress[5]~q ;
wire \dma_1|writeaddress[5]~q ;
wire \dma_2|readaddress[6]~q ;
wire \dma_1|writeaddress[6]~q ;
wire \dma_2|readaddress[7]~q ;
wire \dma_1|writeaddress[7]~q ;
wire \dma_2|readaddress[8]~q ;
wire \dma_1|writeaddress[8]~q ;
wire \dma_2|readaddress[9]~q ;
wire \dma_1|writeaddress[9]~q ;
wire \dma_2|readaddress[10]~q ;
wire \dma_1|writeaddress[10]~q ;
wire \dma_2|readaddress[11]~q ;
wire \dma_1|writeaddress[11]~q ;
wire \dma_2|readaddress[12]~q ;
wire \dma_1|writeaddress[12]~q ;
wire \dma_2|readaddress[13]~q ;
wire \dma_1|writeaddress[13]~q ;
wire \dma_2|readaddress[14]~q ;
wire \dma_1|writeaddress[14]~q ;
wire \dma_1|writeaddress[1]~q ;
wire \dma_1|writeaddress[0]~q ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[1] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[2] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[3] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[4] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[5] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[6] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[7] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[8] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[9] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[10] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[11] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[12] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[13] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[14] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[15] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[16] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[17] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[18] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[19] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[20] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[21] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[22] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[23] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[24] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[25] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[26] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[27] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[28] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[29] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[30] ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[31] ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w0_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w1_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w2_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w3_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w4_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w5_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w6_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w7_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w8_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w9_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w10_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w11_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w12_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w13_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w14_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w15_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w16_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w17_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w18_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w19_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w20_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w21_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w22_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w23_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w24_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w25_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w26_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w27_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w28_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w29_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w30_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w31_n0_mux_dataout~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem_used[7]~q ;
wire \mm_interconnect_1|cmd_mux_001|saved_grant[0]~q ;
wire \dma_1|the_Computer_System_dma_1_mem_read|read_select~q ;
wire \mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|write~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|arvalid~combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|address_taken~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[7]~q ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|fifo_empty~q ;
wire \mm_interconnect_1|cmd_mux|saved_grant[1]~q ;
wire \mm_interconnect_1|cmd_mux|src_valid~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|awvalid~combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|bready~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|data_taken~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|wvalid~combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~0_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~1_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~2_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~3_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~4_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~5_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~6_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~7_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~8_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~9_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~10_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~11_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~12_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~13_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~14_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~15_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~16_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~17_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~18_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~19_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~20_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~21_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~22_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~23_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~24_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~25_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~26_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~27_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~28_combout ;
wire \mm_interconnect_1|cmd_mux_001|src_payload~29_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~0_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~1_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~2_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~3_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~4_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~5_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~6_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~7_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~8_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~9_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~10_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~11_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~12_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~13_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~14_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~15_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~16_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~17_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~18_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~19_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~20_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~21_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~22_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~23_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~24_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~25_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~26_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~27_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~28_combout ;
wire \mm_interconnect_1|cmd_mux|src_payload~29_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_collision~q ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[0]~q ;
wire \dma_2|control[2]~q ;
wire \dma_2|control[0]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~0_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[1]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~1_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[2]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~2_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[3]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~3_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[4]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~4_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[5]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~5_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[6]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~6_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[7]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~7_combout ;
wire \dma_2|write_writedata~0_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[8]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~9_combout ;
wire \dma_2|write_writedata~1_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[9]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~11_combout ;
wire \dma_2|write_writedata~2_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[10]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~13_combout ;
wire \dma_2|write_writedata~3_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[11]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~15_combout ;
wire \dma_2|write_writedata~4_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[12]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~17_combout ;
wire \dma_2|write_writedata~5_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[13]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~19_combout ;
wire \dma_2|write_writedata~6_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[14]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~21_combout ;
wire \dma_2|write_writedata~7_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[15]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~23_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[16]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~25_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[17]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~27_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[18]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~29_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[19]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~31_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[20]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~33_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[21]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~35_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[22]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~37_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[23]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~39_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[24]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~41_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[25]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~43_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[26]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~45_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[27]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~47_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[28]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~49_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[29]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~51_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[30]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~53_combout ;
wire \dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[31]~q ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~55_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~56_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~57_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~58_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~59_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~60_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~61_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~62_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~63_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~64_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~65_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~66_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~67_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~68_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~69_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~70_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~71_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~72_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~73_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~74_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~75_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~76_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~77_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~78_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~79_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~80_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~81_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~82_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~83_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~84_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~85_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~86_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~87_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~1_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~2_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~3_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~4_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~5_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~6_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~7_combout ;
wire \mm_interconnect_0|dma_2_control_port_slave_agent|WideOr0~0_combout ;
wire \mm_interconnect_0|dma_2_control_port_slave_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_agent|WideOr0~0_combout ;
wire \mm_interconnect_0|dma_1_control_port_slave_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_rd_limiter|cmd_sink_ready~1_combout ;
wire \mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[88]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[89]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[90]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[91]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[92]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[93]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[94]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[95]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[96]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[97]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[98]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[99]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~2_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[1]~5_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~8_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~11_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[4]~14_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~17_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~20_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~23_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~26_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~29_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~32_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[11]~35_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~38_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[13]~41_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~44_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[15]~47_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[16]~50_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[17]~53_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[18]~56_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[19]~59_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[20]~62_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[21]~65_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[22]~68_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~71_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[24]~74_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~77_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~80_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~83_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~86_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[29]~89_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~92_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~95_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[88]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[89]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[90]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[91]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[92]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[93]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[94]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[95]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[96]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[97]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[98]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[99]~combout ;
wire \mm_interconnect_2|cmd_mux|saved_grant[0]~q ;
wire \mm_interconnect_2|cmd_mux|saved_grant[1]~q ;
wire \mm_interconnect_2|onchip_sram_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|fifo_empty~q ;
wire \onchip_sram|wren~0_combout ;
wire \rst_controller|r_early_rst~q ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_collision~q ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[0]~q ;
wire \dma_1|control[2]~q ;
wire \dma_1|control[0]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~1_combout ;
wire \mm_interconnect_2|cmd_mux|src_data[38]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[39]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[40]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[41]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[42]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[43]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[44]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[45]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[46]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[47]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[48]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[49]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[50]~combout ;
wire \mm_interconnect_2|cmd_mux|src_data[32]~0_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[1]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~2_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[2]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~3_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[3]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~4_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[4]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~5_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[5]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~6_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[6]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~7_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[7]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~8_combout ;
wire \dma_1|write_writedata~0_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[8]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~9_combout ;
wire \mm_interconnect_2|cmd_mux|src_data[33]~1_combout ;
wire \dma_1|write_writedata~1_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[9]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~10_combout ;
wire \dma_1|write_writedata~2_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[10]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~11_combout ;
wire \dma_1|write_writedata~3_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[11]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~12_combout ;
wire \dma_1|write_writedata~4_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[12]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~13_combout ;
wire \dma_1|write_writedata~5_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[13]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~14_combout ;
wire \dma_1|write_writedata~6_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[14]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~15_combout ;
wire \dma_1|write_writedata~7_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[15]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~16_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[16]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~17_combout ;
wire \mm_interconnect_2|cmd_mux|src_data[34]~2_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[17]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~18_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[18]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~19_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[19]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~20_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[20]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~21_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[21]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~22_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[22]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~23_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[23]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~24_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[24]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~25_combout ;
wire \mm_interconnect_2|cmd_mux|src_data[35]~3_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[25]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~26_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[26]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~27_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[27]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~28_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[28]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~29_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[29]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~30_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[30]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~31_combout ;
wire \dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[31]~q ;
wire \mm_interconnect_2|cmd_mux|src_payload~32_combout ;
wire \rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_1|cmd_mux_001|WideOr1~0_combout ;
wire \rst_controller|r_sync_rst~q ;
wire \dma_1|the_Computer_System_dma_1_mem_read|inc_read~combout ;
wire \mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~0_combout ;
wire \mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~1_combout ;
wire \mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~2_combout ;
wire \mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~3_combout ;
wire \dma_2|the_Computer_System_dma_2_mem_write|fifo_read~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|write_cp_ready~0_combout ;
wire \mm_interconnect_2|rsp_demux|src0_valid~combout ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_agent_rsp_fifo|mem~0_combout ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_agent_rsp_fifo|mem~0_combout ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \onchip_sram|the_altsyncram|auto_generated|address_reg_a[0]~q ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w16_n0_mux_dataout~0_combout ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w17_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w18_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w19_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w20_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w21_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w22_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w23_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w8_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w9_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w10_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w11_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w12_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w13_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w14_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w15_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w24_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w25_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w26_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w27_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w28_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w29_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w30_n0_mux_dataout~0_combout ;
wire \onchip_sram|the_altsyncram|auto_generated|mux4|l1_w31_n0_mux_dataout~0_combout ;
wire \mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \dma_1|dma_ctl_readdata[0]~q ;
wire \dma_2|dma_ctl_readdata[0]~q ;
wire \dma_1|dma_ctl_readdata[1]~q ;
wire \dma_2|dma_ctl_readdata[1]~q ;
wire \dma_1|dma_ctl_readdata[2]~q ;
wire \dma_2|dma_ctl_readdata[2]~q ;
wire \dma_1|dma_ctl_readdata[3]~q ;
wire \dma_2|dma_ctl_readdata[3]~q ;
wire \dma_1|dma_ctl_readdata[4]~q ;
wire \dma_2|dma_ctl_readdata[4]~q ;
wire \dma_1|dma_ctl_readdata[5]~q ;
wire \dma_2|dma_ctl_readdata[5]~q ;
wire \dma_1|dma_ctl_readdata[6]~q ;
wire \dma_2|dma_ctl_readdata[6]~q ;
wire \dma_1|dma_ctl_readdata[7]~q ;
wire \dma_2|dma_ctl_readdata[7]~q ;
wire \dma_1|dma_ctl_readdata[8]~q ;
wire \dma_2|dma_ctl_readdata[8]~q ;
wire \dma_1|dma_ctl_readdata[9]~q ;
wire \dma_2|dma_ctl_readdata[9]~q ;
wire \dma_1|dma_ctl_readdata[10]~q ;
wire \dma_2|dma_ctl_readdata[10]~q ;
wire \dma_1|dma_ctl_readdata[11]~q ;
wire \dma_2|dma_ctl_readdata[11]~q ;
wire \dma_1|dma_ctl_readdata[12]~q ;
wire \dma_2|dma_ctl_readdata[12]~q ;
wire \dma_1|dma_ctl_readdata[13]~q ;
wire \dma_2|dma_ctl_readdata[13]~q ;
wire \dma_1|dma_ctl_readdata[14]~q ;
wire \dma_2|dma_ctl_readdata[14]~q ;
wire \dma_1|dma_ctl_readdata[15]~q ;
wire \dma_2|dma_ctl_readdata[15]~q ;
wire \dma_1|dma_ctl_readdata[16]~q ;
wire \dma_2|dma_ctl_readdata[16]~q ;
wire \dma_1|dma_ctl_readdata[17]~q ;
wire \dma_2|dma_ctl_readdata[17]~q ;
wire \dma_1|dma_ctl_readdata[18]~q ;
wire \dma_2|dma_ctl_readdata[18]~q ;
wire \dma_1|dma_ctl_readdata[19]~q ;
wire \dma_2|dma_ctl_readdata[19]~q ;
wire \dma_1|dma_ctl_readdata[20]~q ;
wire \dma_2|dma_ctl_readdata[20]~q ;
wire \dma_1|dma_ctl_readdata[21]~q ;
wire \dma_2|dma_ctl_readdata[21]~q ;
wire \dma_1|dma_ctl_readdata[22]~q ;
wire \dma_2|dma_ctl_readdata[22]~q ;
wire \dma_1|dma_ctl_readdata[23]~q ;
wire \dma_2|dma_ctl_readdata[23]~q ;
wire \dma_1|dma_ctl_readdata[24]~q ;
wire \dma_2|dma_ctl_readdata[24]~q ;
wire \dma_1|dma_ctl_readdata[25]~q ;
wire \dma_2|dma_ctl_readdata[25]~q ;
wire \dma_1|dma_ctl_readdata[26]~q ;
wire \dma_2|dma_ctl_readdata[26]~q ;
wire \dma_1|dma_ctl_readdata[27]~q ;
wire \dma_2|dma_ctl_readdata[27]~q ;
wire \dma_1|dma_ctl_readdata[28]~q ;
wire \dma_2|dma_ctl_readdata[28]~q ;
wire \dma_1|dma_ctl_readdata[29]~q ;
wire \dma_2|dma_ctl_readdata[29]~q ;
wire \dma_1|dma_ctl_readdata[30]~q ;
wire \dma_2|dma_ctl_readdata[30]~q ;
wire \dma_1|dma_ctl_readdata[31]~q ;
wire \dma_2|dma_ctl_readdata[31]~q ;
wire \dma_2|the_Computer_System_dma_2_mem_read|read_select~q ;
wire \mm_interconnect_2|onchip_sram_s1_translator|read_latency_shift_reg~0_combout ;
wire \mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~4_combout ;
wire \mm_interconnect_1|rsp_demux|src0_valid~1_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[8]~0_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[8]~1_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[16]~4_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[24]~7_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[0]~8_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[0]~9_combout ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_1|rsp_mux|src_data[9]~10_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[9]~11_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[17]~14_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[25]~17_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[1]~18_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[1]~19_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[10]~20_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[10]~21_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[18]~24_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[26]~27_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[2]~28_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[2]~29_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[11]~30_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[11]~31_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[19]~34_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[27]~37_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[3]~38_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[3]~39_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[12]~40_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[12]~41_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[20]~44_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[28]~47_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[4]~48_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[4]~49_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[13]~50_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[13]~51_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[21]~54_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[29]~57_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[5]~58_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[5]~59_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[14]~60_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[14]~61_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[22]~64_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[30]~67_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[6]~68_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[6]~69_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[15]~70_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[15]~71_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[23]~74_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[31]~77_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[7]~78_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[7]~79_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[8]~80_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[9]~81_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[10]~82_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[11]~83_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[12]~84_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[13]~85_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[14]~86_combout ;
wire \mm_interconnect_1|rsp_mux|src_data[15]~87_combout ;
wire \mm_interconnect_2|cmd_mux|src_data[51]~combout ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;
wire \arm_a9_hps|hps_io|border|intermediate[0] ;
wire \arm_a9_hps|hps_io|border|intermediate[1] ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;
wire \arm_a9_hps|hps_io|border|emac1_inst~emac_phy_txd ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;
wire \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SCLK ;
wire \arm_a9_hps|hps_io|border|intermediate[2] ;
wire \arm_a9_hps|hps_io|border|intermediate[4] ;
wire \arm_a9_hps|hps_io|border|intermediate[6] ;
wire \arm_a9_hps|hps_io|border|intermediate[8] ;
wire \arm_a9_hps|hps_io|border|intermediate[3] ;
wire \arm_a9_hps|hps_io|border|intermediate[5] ;
wire \arm_a9_hps|hps_io|border|intermediate[7] ;
wire \arm_a9_hps|hps_io|border|intermediate[9] ;
wire \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;
wire \arm_a9_hps|hps_io|border|sdio_inst~sdmmc_cclk ;
wire \arm_a9_hps|hps_io|border|intermediate[10] ;
wire \arm_a9_hps|hps_io|border|intermediate[11] ;
wire \arm_a9_hps|hps_io|border|intermediate[12] ;
wire \arm_a9_hps|hps_io|border|intermediate[14] ;
wire \arm_a9_hps|hps_io|border|intermediate[16] ;
wire \arm_a9_hps|hps_io|border|intermediate[18] ;
wire \arm_a9_hps|hps_io|border|intermediate[13] ;
wire \arm_a9_hps|hps_io|border|intermediate[15] ;
wire \arm_a9_hps|hps_io|border|intermediate[17] ;
wire \arm_a9_hps|hps_io|border|intermediate[19] ;
wire \arm_a9_hps|hps_io|border|usb1_inst~usb_ulpi_stp ;
wire \arm_a9_hps|hps_io|border|intermediate[20] ;
wire \arm_a9_hps|hps_io|border|intermediate[22] ;
wire \arm_a9_hps|hps_io|border|intermediate[24] ;
wire \arm_a9_hps|hps_io|border|intermediate[26] ;
wire \arm_a9_hps|hps_io|border|intermediate[28] ;
wire \arm_a9_hps|hps_io|border|intermediate[30] ;
wire \arm_a9_hps|hps_io|border|intermediate[32] ;
wire \arm_a9_hps|hps_io|border|intermediate[34] ;
wire \arm_a9_hps|hps_io|border|intermediate[21] ;
wire \arm_a9_hps|hps_io|border|intermediate[23] ;
wire \arm_a9_hps|hps_io|border|intermediate[25] ;
wire \arm_a9_hps|hps_io|border|intermediate[27] ;
wire \arm_a9_hps|hps_io|border|intermediate[29] ;
wire \arm_a9_hps|hps_io|border|intermediate[31] ;
wire \arm_a9_hps|hps_io|border|intermediate[33] ;
wire \arm_a9_hps|hps_io|border|intermediate[35] ;
wire \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;
wire \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;
wire \arm_a9_hps|hps_io|border|intermediate[36] ;
wire \arm_a9_hps|hps_io|border|intermediate[37] ;
wire \arm_a9_hps|hps_io|border|uart0_inst~uart_txd ;
wire \arm_a9_hps|hps_io|border|intermediate[39] ;
wire \arm_a9_hps|hps_io|border|intermediate[38] ;
wire \arm_a9_hps|hps_io|border|intermediate[41] ;
wire \arm_a9_hps|hps_io|border|intermediate[40] ;
wire \arm_a9_hps|hps_io|border|intermediate[42] ;
wire \arm_a9_hps|hps_io|border|intermediate[43] ;
wire \arm_a9_hps|hps_io|border|intermediate[44] ;
wire \arm_a9_hps|hps_io|border|intermediate[46] ;
wire \arm_a9_hps|hps_io|border|intermediate[48] ;
wire \arm_a9_hps|hps_io|border|intermediate[50] ;
wire \arm_a9_hps|hps_io|border|intermediate[52] ;
wire \arm_a9_hps|hps_io|border|intermediate[54] ;
wire \arm_a9_hps|hps_io|border|intermediate[45] ;
wire \arm_a9_hps|hps_io|border|intermediate[47] ;
wire \arm_a9_hps|hps_io|border|intermediate[49] ;
wire \arm_a9_hps|hps_io|border|intermediate[51] ;
wire \arm_a9_hps|hps_io|border|intermediate[53] ;
wire \arm_a9_hps|hps_io|border|intermediate[55] ;
wire \arm_a9_hps|hps_io|border|intermediate[56] ;
wire \arm_a9_hps|hps_io|border|intermediate[57] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \onchip_sram_reset2_reset~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o ;
wire \hps_f2h_irq0_irq[0]~input_o ;
wire \hps_f2h_irq0_irq[1]~input_o ;
wire \hps_f2h_irq0_irq[2]~input_o ;
wire \hps_f2h_irq0_irq[3]~input_o ;
wire \hps_f2h_irq0_irq[4]~input_o ;
wire \hps_f2h_irq0_irq[5]~input_o ;
wire \hps_f2h_irq0_irq[6]~input_o ;
wire \hps_f2h_irq0_irq[7]~input_o ;
wire \hps_f2h_irq0_irq[8]~input_o ;
wire \hps_f2h_irq0_irq[9]~input_o ;
wire \hps_f2h_irq0_irq[10]~input_o ;
wire \hps_f2h_irq0_irq[11]~input_o ;
wire \hps_f2h_irq0_irq[12]~input_o ;
wire \hps_f2h_irq0_irq[13]~input_o ;
wire \hps_f2h_irq0_irq[14]~input_o ;
wire \hps_f2h_irq0_irq[15]~input_o ;
wire \hps_f2h_irq0_irq[16]~input_o ;
wire \hps_f2h_irq0_irq[17]~input_o ;
wire \hps_f2h_irq0_irq[18]~input_o ;
wire \hps_f2h_irq0_irq[19]~input_o ;
wire \hps_f2h_irq0_irq[20]~input_o ;
wire \hps_f2h_irq0_irq[21]~input_o ;
wire \hps_f2h_irq0_irq[22]~input_o ;
wire \hps_f2h_irq0_irq[23]~input_o ;
wire \hps_f2h_irq0_irq[24]~input_o ;
wire \hps_f2h_irq0_irq[25]~input_o ;
wire \hps_f2h_irq0_irq[26]~input_o ;
wire \hps_f2h_irq0_irq[27]~input_o ;
wire \hps_f2h_irq0_irq[28]~input_o ;
wire \hps_f2h_irq0_irq[29]~input_o ;
wire \hps_f2h_irq0_irq[30]~input_o ;
wire \hps_f2h_irq0_irq[31]~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD0~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD1~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD2~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD3~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CLK~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CTL~input_o ;
wire \hps_io_hps_io_spim1_inst_MISO~input_o ;
wire \hps_io_hps_io_uart0_inst_RX~input_o ;
wire \hps_io_hps_io_usb1_inst_CLK~input_o ;
wire \hps_io_hps_io_usb1_inst_DIR~input_o ;
wire \hps_io_hps_io_usb1_inst_NXT~input_o ;
wire \memory_oct_rzqin~input_o ;
wire \onchip_sram_s2_address[13]~input_o ;
wire \onchip_sram_s2_chipselect~input_o ;
wire \onchip_sram_s2_write~input_o ;
wire \onchip_sram_clk2_clk~input_o ;
wire \onchip_sram_reset2_reset_req~input_o ;
wire \onchip_sram_s2_clken~input_o ;
wire \onchip_sram_s2_writedata[0]~input_o ;
wire \onchip_sram_s2_address[0]~input_o ;
wire \onchip_sram_s2_address[1]~input_o ;
wire \onchip_sram_s2_address[2]~input_o ;
wire \onchip_sram_s2_address[3]~input_o ;
wire \onchip_sram_s2_address[4]~input_o ;
wire \onchip_sram_s2_address[5]~input_o ;
wire \onchip_sram_s2_address[6]~input_o ;
wire \onchip_sram_s2_address[7]~input_o ;
wire \onchip_sram_s2_address[8]~input_o ;
wire \onchip_sram_s2_address[9]~input_o ;
wire \onchip_sram_s2_address[10]~input_o ;
wire \onchip_sram_s2_address[11]~input_o ;
wire \onchip_sram_s2_address[12]~input_o ;
wire \onchip_sram_s2_byteenable[0]~input_o ;
wire \onchip_sram_s2_writedata[1]~input_o ;
wire \onchip_sram_s2_writedata[2]~input_o ;
wire \onchip_sram_s2_writedata[3]~input_o ;
wire \onchip_sram_s2_writedata[4]~input_o ;
wire \onchip_sram_s2_writedata[5]~input_o ;
wire \onchip_sram_s2_writedata[6]~input_o ;
wire \onchip_sram_s2_writedata[7]~input_o ;
wire \onchip_sram_s2_writedata[8]~input_o ;
wire \onchip_sram_s2_byteenable[1]~input_o ;
wire \onchip_sram_s2_writedata[9]~input_o ;
wire \onchip_sram_s2_writedata[10]~input_o ;
wire \onchip_sram_s2_writedata[11]~input_o ;
wire \onchip_sram_s2_writedata[12]~input_o ;
wire \onchip_sram_s2_writedata[13]~input_o ;
wire \onchip_sram_s2_writedata[14]~input_o ;
wire \onchip_sram_s2_writedata[15]~input_o ;
wire \onchip_sram_s2_writedata[16]~input_o ;
wire \onchip_sram_s2_byteenable[2]~input_o ;
wire \onchip_sram_s2_writedata[17]~input_o ;
wire \onchip_sram_s2_writedata[18]~input_o ;
wire \onchip_sram_s2_writedata[19]~input_o ;
wire \onchip_sram_s2_writedata[20]~input_o ;
wire \onchip_sram_s2_writedata[21]~input_o ;
wire \onchip_sram_s2_writedata[22]~input_o ;
wire \onchip_sram_s2_writedata[23]~input_o ;
wire \onchip_sram_s2_writedata[24]~input_o ;
wire \onchip_sram_s2_byteenable[3]~input_o ;
wire \onchip_sram_s2_writedata[25]~input_o ;
wire \onchip_sram_s2_writedata[26]~input_o ;
wire \onchip_sram_s2_writedata[27]~input_o ;
wire \onchip_sram_s2_writedata[28]~input_o ;
wire \onchip_sram_s2_writedata[29]~input_o ;
wire \onchip_sram_s2_writedata[30]~input_o ;
wire \onchip_sram_s2_writedata[31]~input_o ;
wire \system_pll_ref_clk_clk~input_o ;
wire \system_pll_ref_reset_reset~input_o ;


Computer_System_Computer_System_ARM_A9_HPS arm_a9_hps(
	.h2f_rst_n_0(\arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ),
	.f2h_ARREADY_0(\arm_a9_hps|fpga_interfaces|f2h_ARREADY[0] ),
	.f2h_AWREADY_0(\arm_a9_hps|fpga_interfaces|f2h_AWREADY[0] ),
	.f2h_BVALID_0(\arm_a9_hps|fpga_interfaces|f2h_BVALID[0] ),
	.f2h_RVALID_0(\arm_a9_hps|fpga_interfaces|f2h_RVALID[0] ),
	.f2h_WREADY_0(\arm_a9_hps|fpga_interfaces|f2h_WREADY[0] ),
	.f2h_RDATA_0(\arm_a9_hps|fpga_interfaces|f2h_RDATA[0] ),
	.f2h_RDATA_1(\arm_a9_hps|fpga_interfaces|f2h_RDATA[1] ),
	.f2h_RDATA_2(\arm_a9_hps|fpga_interfaces|f2h_RDATA[2] ),
	.f2h_RDATA_3(\arm_a9_hps|fpga_interfaces|f2h_RDATA[3] ),
	.f2h_RDATA_4(\arm_a9_hps|fpga_interfaces|f2h_RDATA[4] ),
	.f2h_RDATA_5(\arm_a9_hps|fpga_interfaces|f2h_RDATA[5] ),
	.f2h_RDATA_6(\arm_a9_hps|fpga_interfaces|f2h_RDATA[6] ),
	.f2h_RDATA_7(\arm_a9_hps|fpga_interfaces|f2h_RDATA[7] ),
	.f2h_RDATA_8(\arm_a9_hps|fpga_interfaces|f2h_RDATA[8] ),
	.f2h_RDATA_9(\arm_a9_hps|fpga_interfaces|f2h_RDATA[9] ),
	.f2h_RDATA_10(\arm_a9_hps|fpga_interfaces|f2h_RDATA[10] ),
	.f2h_RDATA_11(\arm_a9_hps|fpga_interfaces|f2h_RDATA[11] ),
	.f2h_RDATA_12(\arm_a9_hps|fpga_interfaces|f2h_RDATA[12] ),
	.f2h_RDATA_13(\arm_a9_hps|fpga_interfaces|f2h_RDATA[13] ),
	.f2h_RDATA_14(\arm_a9_hps|fpga_interfaces|f2h_RDATA[14] ),
	.f2h_RDATA_15(\arm_a9_hps|fpga_interfaces|f2h_RDATA[15] ),
	.f2h_RDATA_16(\arm_a9_hps|fpga_interfaces|f2h_RDATA[16] ),
	.f2h_RDATA_17(\arm_a9_hps|fpga_interfaces|f2h_RDATA[17] ),
	.f2h_RDATA_18(\arm_a9_hps|fpga_interfaces|f2h_RDATA[18] ),
	.f2h_RDATA_19(\arm_a9_hps|fpga_interfaces|f2h_RDATA[19] ),
	.f2h_RDATA_20(\arm_a9_hps|fpga_interfaces|f2h_RDATA[20] ),
	.f2h_RDATA_21(\arm_a9_hps|fpga_interfaces|f2h_RDATA[21] ),
	.f2h_RDATA_22(\arm_a9_hps|fpga_interfaces|f2h_RDATA[22] ),
	.f2h_RDATA_23(\arm_a9_hps|fpga_interfaces|f2h_RDATA[23] ),
	.f2h_RDATA_24(\arm_a9_hps|fpga_interfaces|f2h_RDATA[24] ),
	.f2h_RDATA_25(\arm_a9_hps|fpga_interfaces|f2h_RDATA[25] ),
	.f2h_RDATA_26(\arm_a9_hps|fpga_interfaces|f2h_RDATA[26] ),
	.f2h_RDATA_27(\arm_a9_hps|fpga_interfaces|f2h_RDATA[27] ),
	.f2h_RDATA_28(\arm_a9_hps|fpga_interfaces|f2h_RDATA[28] ),
	.f2h_RDATA_29(\arm_a9_hps|fpga_interfaces|f2h_RDATA[29] ),
	.f2h_RDATA_30(\arm_a9_hps|fpga_interfaces|f2h_RDATA[30] ),
	.f2h_RDATA_31(\arm_a9_hps|fpga_interfaces|f2h_RDATA[31] ),
	.f2h_RDATA_32(\arm_a9_hps|fpga_interfaces|f2h_RDATA[32] ),
	.f2h_RDATA_33(\arm_a9_hps|fpga_interfaces|f2h_RDATA[33] ),
	.f2h_RDATA_34(\arm_a9_hps|fpga_interfaces|f2h_RDATA[34] ),
	.f2h_RDATA_35(\arm_a9_hps|fpga_interfaces|f2h_RDATA[35] ),
	.f2h_RDATA_36(\arm_a9_hps|fpga_interfaces|f2h_RDATA[36] ),
	.f2h_RDATA_37(\arm_a9_hps|fpga_interfaces|f2h_RDATA[37] ),
	.f2h_RDATA_38(\arm_a9_hps|fpga_interfaces|f2h_RDATA[38] ),
	.f2h_RDATA_39(\arm_a9_hps|fpga_interfaces|f2h_RDATA[39] ),
	.f2h_RDATA_40(\arm_a9_hps|fpga_interfaces|f2h_RDATA[40] ),
	.f2h_RDATA_41(\arm_a9_hps|fpga_interfaces|f2h_RDATA[41] ),
	.f2h_RDATA_42(\arm_a9_hps|fpga_interfaces|f2h_RDATA[42] ),
	.f2h_RDATA_43(\arm_a9_hps|fpga_interfaces|f2h_RDATA[43] ),
	.f2h_RDATA_44(\arm_a9_hps|fpga_interfaces|f2h_RDATA[44] ),
	.f2h_RDATA_45(\arm_a9_hps|fpga_interfaces|f2h_RDATA[45] ),
	.f2h_RDATA_46(\arm_a9_hps|fpga_interfaces|f2h_RDATA[46] ),
	.f2h_RDATA_47(\arm_a9_hps|fpga_interfaces|f2h_RDATA[47] ),
	.f2h_RDATA_48(\arm_a9_hps|fpga_interfaces|f2h_RDATA[48] ),
	.f2h_RDATA_49(\arm_a9_hps|fpga_interfaces|f2h_RDATA[49] ),
	.f2h_RDATA_50(\arm_a9_hps|fpga_interfaces|f2h_RDATA[50] ),
	.f2h_RDATA_51(\arm_a9_hps|fpga_interfaces|f2h_RDATA[51] ),
	.f2h_RDATA_52(\arm_a9_hps|fpga_interfaces|f2h_RDATA[52] ),
	.f2h_RDATA_53(\arm_a9_hps|fpga_interfaces|f2h_RDATA[53] ),
	.f2h_RDATA_54(\arm_a9_hps|fpga_interfaces|f2h_RDATA[54] ),
	.f2h_RDATA_55(\arm_a9_hps|fpga_interfaces|f2h_RDATA[55] ),
	.f2h_RDATA_56(\arm_a9_hps|fpga_interfaces|f2h_RDATA[56] ),
	.f2h_RDATA_57(\arm_a9_hps|fpga_interfaces|f2h_RDATA[57] ),
	.f2h_RDATA_58(\arm_a9_hps|fpga_interfaces|f2h_RDATA[58] ),
	.f2h_RDATA_59(\arm_a9_hps|fpga_interfaces|f2h_RDATA[59] ),
	.f2h_RDATA_60(\arm_a9_hps|fpga_interfaces|f2h_RDATA[60] ),
	.f2h_RDATA_61(\arm_a9_hps|fpga_interfaces|f2h_RDATA[61] ),
	.f2h_RDATA_62(\arm_a9_hps|fpga_interfaces|f2h_RDATA[62] ),
	.f2h_RDATA_63(\arm_a9_hps|fpga_interfaces|f2h_RDATA[63] ),
	.h2f_lw_ARVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARADDR_5(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[5] ),
	.h2f_lw_ARBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWADDR_5(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[5] ),
	.h2f_lw_AWBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.saved_grant_0(\mm_interconnect_1|cmd_mux_001|saved_grant[0]~q ),
	.arvalid(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|arvalid~combout ),
	.saved_grant_1(\mm_interconnect_1|cmd_mux|saved_grant[1]~q ),
	.awvalid(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|awvalid~combout ),
	.bready(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|bready~0_combout ),
	.wvalid(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|wvalid~combout ),
	.src_payload(\mm_interconnect_1|cmd_mux_001|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_1|cmd_mux_001|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_1|cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_1|cmd_mux_001|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_1|cmd_mux_001|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_1|cmd_mux_001|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_1|cmd_mux_001|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_1|cmd_mux_001|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_1|cmd_mux_001|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_1|cmd_mux_001|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_1|cmd_mux_001|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_1|cmd_mux_001|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_1|cmd_mux_001|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_1|cmd_mux_001|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_1|cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_1|cmd_mux_001|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_1|cmd_mux_001|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_1|cmd_mux_001|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_1|cmd_mux_001|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_1|cmd_mux_001|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_1|cmd_mux_001|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_1|cmd_mux_001|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_1|cmd_mux_001|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_1|cmd_mux_001|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_1|cmd_mux_001|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_1|cmd_mux_001|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_1|cmd_mux_001|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_1|cmd_mux_001|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_1|cmd_mux_001|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_1|cmd_mux_001|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_1|cmd_mux|src_payload~0_combout ),
	.src_payload31(\mm_interconnect_1|cmd_mux|src_payload~1_combout ),
	.src_payload32(\mm_interconnect_1|cmd_mux|src_payload~2_combout ),
	.src_payload33(\mm_interconnect_1|cmd_mux|src_payload~3_combout ),
	.src_payload34(\mm_interconnect_1|cmd_mux|src_payload~4_combout ),
	.src_payload35(\mm_interconnect_1|cmd_mux|src_payload~5_combout ),
	.src_payload36(\mm_interconnect_1|cmd_mux|src_payload~6_combout ),
	.src_payload37(\mm_interconnect_1|cmd_mux|src_payload~7_combout ),
	.src_payload38(\mm_interconnect_1|cmd_mux|src_payload~8_combout ),
	.src_payload39(\mm_interconnect_1|cmd_mux|src_payload~9_combout ),
	.src_payload40(\mm_interconnect_1|cmd_mux|src_payload~10_combout ),
	.src_payload41(\mm_interconnect_1|cmd_mux|src_payload~11_combout ),
	.src_payload42(\mm_interconnect_1|cmd_mux|src_payload~12_combout ),
	.src_payload43(\mm_interconnect_1|cmd_mux|src_payload~13_combout ),
	.src_payload44(\mm_interconnect_1|cmd_mux|src_payload~14_combout ),
	.src_payload45(\mm_interconnect_1|cmd_mux|src_payload~15_combout ),
	.src_payload46(\mm_interconnect_1|cmd_mux|src_payload~16_combout ),
	.src_payload47(\mm_interconnect_1|cmd_mux|src_payload~17_combout ),
	.src_payload48(\mm_interconnect_1|cmd_mux|src_payload~18_combout ),
	.src_payload49(\mm_interconnect_1|cmd_mux|src_payload~19_combout ),
	.src_payload50(\mm_interconnect_1|cmd_mux|src_payload~20_combout ),
	.src_payload51(\mm_interconnect_1|cmd_mux|src_payload~21_combout ),
	.src_payload52(\mm_interconnect_1|cmd_mux|src_payload~22_combout ),
	.src_payload53(\mm_interconnect_1|cmd_mux|src_payload~23_combout ),
	.src_payload54(\mm_interconnect_1|cmd_mux|src_payload~24_combout ),
	.src_payload55(\mm_interconnect_1|cmd_mux|src_payload~25_combout ),
	.src_payload56(\mm_interconnect_1|cmd_mux|src_payload~26_combout ),
	.src_payload57(\mm_interconnect_1|cmd_mux|src_payload~27_combout ),
	.src_payload58(\mm_interconnect_1|cmd_mux|src_payload~28_combout ),
	.src_payload59(\mm_interconnect_1|cmd_mux|src_payload~29_combout ),
	.ShiftLeft1(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~0_combout ),
	.ShiftLeft11(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~1_combout ),
	.ShiftLeft12(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~2_combout ),
	.ShiftLeft13(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~3_combout ),
	.ShiftLeft14(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~4_combout ),
	.ShiftLeft15(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~5_combout ),
	.ShiftLeft16(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~6_combout ),
	.ShiftLeft17(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~7_combout ),
	.ShiftLeft18(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~9_combout ),
	.ShiftLeft19(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~11_combout ),
	.ShiftLeft110(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~13_combout ),
	.ShiftLeft111(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~15_combout ),
	.ShiftLeft112(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~17_combout ),
	.ShiftLeft113(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~19_combout ),
	.ShiftLeft114(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~21_combout ),
	.ShiftLeft115(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~23_combout ),
	.ShiftLeft116(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~25_combout ),
	.ShiftLeft117(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~27_combout ),
	.ShiftLeft118(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~29_combout ),
	.ShiftLeft119(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~31_combout ),
	.ShiftLeft120(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~33_combout ),
	.ShiftLeft121(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~35_combout ),
	.ShiftLeft122(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~37_combout ),
	.ShiftLeft123(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~39_combout ),
	.ShiftLeft124(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~41_combout ),
	.ShiftLeft125(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~43_combout ),
	.ShiftLeft126(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~45_combout ),
	.ShiftLeft127(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~47_combout ),
	.ShiftLeft128(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~49_combout ),
	.ShiftLeft129(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~51_combout ),
	.ShiftLeft130(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~53_combout ),
	.ShiftLeft131(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~55_combout ),
	.ShiftLeft132(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~56_combout ),
	.ShiftLeft133(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~57_combout ),
	.ShiftLeft134(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~58_combout ),
	.ShiftLeft135(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~59_combout ),
	.ShiftLeft136(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~60_combout ),
	.ShiftLeft137(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~61_combout ),
	.ShiftLeft138(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~62_combout ),
	.ShiftLeft139(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~63_combout ),
	.ShiftLeft140(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~64_combout ),
	.ShiftLeft141(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~65_combout ),
	.ShiftLeft142(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~66_combout ),
	.ShiftLeft143(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~67_combout ),
	.ShiftLeft144(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~68_combout ),
	.ShiftLeft145(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~69_combout ),
	.ShiftLeft146(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~70_combout ),
	.ShiftLeft147(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~71_combout ),
	.ShiftLeft148(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~72_combout ),
	.ShiftLeft149(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~73_combout ),
	.ShiftLeft150(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~74_combout ),
	.ShiftLeft151(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~75_combout ),
	.ShiftLeft152(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~76_combout ),
	.ShiftLeft153(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~77_combout ),
	.ShiftLeft154(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~78_combout ),
	.ShiftLeft155(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~79_combout ),
	.ShiftLeft156(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~80_combout ),
	.ShiftLeft157(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~81_combout ),
	.ShiftLeft158(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~82_combout ),
	.ShiftLeft159(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~83_combout ),
	.ShiftLeft160(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~84_combout ),
	.ShiftLeft161(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~85_combout ),
	.ShiftLeft162(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~86_combout ),
	.ShiftLeft163(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~87_combout ),
	.ShiftLeft0(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~0_combout ),
	.ShiftLeft01(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~1_combout ),
	.ShiftLeft02(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~2_combout ),
	.ShiftLeft03(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~3_combout ),
	.ShiftLeft04(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~4_combout ),
	.ShiftLeft05(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~5_combout ),
	.ShiftLeft06(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~6_combout ),
	.ShiftLeft07(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~7_combout ),
	.cmd_sink_ready(\mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_rd_limiter|cmd_sink_ready~1_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.nonposted_cmd_accepted1(\mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ),
	.src_data_88(\mm_interconnect_0|rsp_mux|src_data[88]~combout ),
	.src_data_89(\mm_interconnect_0|rsp_mux|src_data[89]~combout ),
	.src_data_90(\mm_interconnect_0|rsp_mux|src_data[90]~combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux|src_data[91]~combout ),
	.src_data_92(\mm_interconnect_0|rsp_mux|src_data[92]~combout ),
	.src_data_93(\mm_interconnect_0|rsp_mux|src_data[93]~combout ),
	.src_data_94(\mm_interconnect_0|rsp_mux|src_data[94]~combout ),
	.src_data_95(\mm_interconnect_0|rsp_mux|src_data[95]~combout ),
	.src_data_96(\mm_interconnect_0|rsp_mux|src_data[96]~combout ),
	.src_data_97(\mm_interconnect_0|rsp_mux|src_data[97]~combout ),
	.src_data_98(\mm_interconnect_0|rsp_mux|src_data[98]~combout ),
	.src_data_99(\mm_interconnect_0|rsp_mux|src_data[99]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~2_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux_001|src_data[1]~5_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~8_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux_001|src_data[3]~11_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux_001|src_data[4]~14_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~17_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~20_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~23_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~26_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~29_combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~32_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[11]~35_combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~38_combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux_001|src_data[13]~41_combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~44_combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~47_combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~50_combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~53_combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~56_combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~59_combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux_001|src_data[20]~62_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[21]~65_combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~68_combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~71_combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~74_combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~77_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~80_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~83_combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~86_combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~89_combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~92_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[31]~95_combout ),
	.src_data_881(\mm_interconnect_0|rsp_mux_001|src_data[88]~combout ),
	.src_data_891(\mm_interconnect_0|rsp_mux_001|src_data[89]~combout ),
	.src_data_901(\mm_interconnect_0|rsp_mux_001|src_data[90]~combout ),
	.src_data_911(\mm_interconnect_0|rsp_mux_001|src_data[91]~combout ),
	.src_data_921(\mm_interconnect_0|rsp_mux_001|src_data[92]~combout ),
	.src_data_931(\mm_interconnect_0|rsp_mux_001|src_data[93]~combout ),
	.src_data_941(\mm_interconnect_0|rsp_mux_001|src_data[94]~combout ),
	.src_data_951(\mm_interconnect_0|rsp_mux_001|src_data[95]~combout ),
	.src_data_961(\mm_interconnect_0|rsp_mux_001|src_data[96]~combout ),
	.src_data_971(\mm_interconnect_0|rsp_mux_001|src_data[97]~combout ),
	.src_data_981(\mm_interconnect_0|rsp_mux_001|src_data[98]~combout ),
	.src_data_991(\mm_interconnect_0|rsp_mux_001|src_data[99]~combout ),
	.emac1_inst(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ),
	.emac1_inst1(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ),
	.intermediate_0(\arm_a9_hps|hps_io|border|intermediate[0] ),
	.intermediate_1(\arm_a9_hps|hps_io|border|intermediate[1] ),
	.emac1_inst2(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ),
	.emac1_inst3(\arm_a9_hps|hps_io|border|emac1_inst~emac_phy_txd ),
	.emac1_inst4(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ),
	.emac1_inst5(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ),
	.emac1_inst6(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ),
	.qspi_inst(\arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SCLK ),
	.intermediate_2(\arm_a9_hps|hps_io|border|intermediate[2] ),
	.intermediate_4(\arm_a9_hps|hps_io|border|intermediate[4] ),
	.intermediate_6(\arm_a9_hps|hps_io|border|intermediate[6] ),
	.intermediate_8(\arm_a9_hps|hps_io|border|intermediate[8] ),
	.intermediate_3(\arm_a9_hps|hps_io|border|intermediate[3] ),
	.intermediate_5(\arm_a9_hps|hps_io|border|intermediate[5] ),
	.intermediate_7(\arm_a9_hps|hps_io|border|intermediate[7] ),
	.intermediate_9(\arm_a9_hps|hps_io|border|intermediate[9] ),
	.qspi_inst1(\arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SS_N0 ),
	.sdio_inst(\arm_a9_hps|hps_io|border|sdio_inst~sdmmc_cclk ),
	.intermediate_10(\arm_a9_hps|hps_io|border|intermediate[10] ),
	.intermediate_11(\arm_a9_hps|hps_io|border|intermediate[11] ),
	.intermediate_12(\arm_a9_hps|hps_io|border|intermediate[12] ),
	.intermediate_14(\arm_a9_hps|hps_io|border|intermediate[14] ),
	.intermediate_16(\arm_a9_hps|hps_io|border|intermediate[16] ),
	.intermediate_18(\arm_a9_hps|hps_io|border|intermediate[18] ),
	.intermediate_13(\arm_a9_hps|hps_io|border|intermediate[13] ),
	.intermediate_15(\arm_a9_hps|hps_io|border|intermediate[15] ),
	.intermediate_17(\arm_a9_hps|hps_io|border|intermediate[17] ),
	.intermediate_19(\arm_a9_hps|hps_io|border|intermediate[19] ),
	.usb1_inst(\arm_a9_hps|hps_io|border|usb1_inst~usb_ulpi_stp ),
	.intermediate_20(\arm_a9_hps|hps_io|border|intermediate[20] ),
	.intermediate_22(\arm_a9_hps|hps_io|border|intermediate[22] ),
	.intermediate_24(\arm_a9_hps|hps_io|border|intermediate[24] ),
	.intermediate_26(\arm_a9_hps|hps_io|border|intermediate[26] ),
	.intermediate_28(\arm_a9_hps|hps_io|border|intermediate[28] ),
	.intermediate_30(\arm_a9_hps|hps_io|border|intermediate[30] ),
	.intermediate_32(\arm_a9_hps|hps_io|border|intermediate[32] ),
	.intermediate_34(\arm_a9_hps|hps_io|border|intermediate[34] ),
	.intermediate_21(\arm_a9_hps|hps_io|border|intermediate[21] ),
	.intermediate_23(\arm_a9_hps|hps_io|border|intermediate[23] ),
	.intermediate_25(\arm_a9_hps|hps_io|border|intermediate[25] ),
	.intermediate_27(\arm_a9_hps|hps_io|border|intermediate[27] ),
	.intermediate_29(\arm_a9_hps|hps_io|border|intermediate[29] ),
	.intermediate_31(\arm_a9_hps|hps_io|border|intermediate[31] ),
	.intermediate_33(\arm_a9_hps|hps_io|border|intermediate[33] ),
	.intermediate_35(\arm_a9_hps|hps_io|border|intermediate[35] ),
	.spim1_inst(\arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ),
	.spim1_inst1(\arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ),
	.intermediate_36(\arm_a9_hps|hps_io|border|intermediate[36] ),
	.intermediate_37(\arm_a9_hps|hps_io|border|intermediate[37] ),
	.uart0_inst(\arm_a9_hps|hps_io|border|uart0_inst~uart_txd ),
	.intermediate_39(\arm_a9_hps|hps_io|border|intermediate[39] ),
	.intermediate_38(\arm_a9_hps|hps_io|border|intermediate[38] ),
	.intermediate_41(\arm_a9_hps|hps_io|border|intermediate[41] ),
	.intermediate_40(\arm_a9_hps|hps_io|border|intermediate[40] ),
	.intermediate_42(\arm_a9_hps|hps_io|border|intermediate[42] ),
	.intermediate_43(\arm_a9_hps|hps_io|border|intermediate[43] ),
	.intermediate_44(\arm_a9_hps|hps_io|border|intermediate[44] ),
	.intermediate_46(\arm_a9_hps|hps_io|border|intermediate[46] ),
	.intermediate_48(\arm_a9_hps|hps_io|border|intermediate[48] ),
	.intermediate_50(\arm_a9_hps|hps_io|border|intermediate[50] ),
	.intermediate_52(\arm_a9_hps|hps_io|border|intermediate[52] ),
	.intermediate_54(\arm_a9_hps|hps_io|border|intermediate[54] ),
	.intermediate_45(\arm_a9_hps|hps_io|border|intermediate[45] ),
	.intermediate_47(\arm_a9_hps|hps_io|border|intermediate[47] ),
	.intermediate_49(\arm_a9_hps|hps_io|border|intermediate[49] ),
	.intermediate_51(\arm_a9_hps|hps_io|border|intermediate[51] ),
	.intermediate_53(\arm_a9_hps|hps_io|border|intermediate[53] ),
	.intermediate_55(\arm_a9_hps|hps_io|border|intermediate[55] ),
	.intermediate_56(\arm_a9_hps|hps_io|border|intermediate[56] ),
	.intermediate_57(\arm_a9_hps|hps_io|border|intermediate[57] ),
	.parallelterminationcontrol_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ),
	.parallelterminationcontrol_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ),
	.parallelterminationcontrol_2(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ),
	.parallelterminationcontrol_3(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ),
	.parallelterminationcontrol_4(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ),
	.parallelterminationcontrol_5(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ),
	.parallelterminationcontrol_6(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ),
	.parallelterminationcontrol_7(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ),
	.parallelterminationcontrol_8(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ),
	.parallelterminationcontrol_9(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ),
	.parallelterminationcontrol_10(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ),
	.parallelterminationcontrol_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ),
	.parallelterminationcontrol_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ),
	.parallelterminationcontrol_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ),
	.parallelterminationcontrol_14(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ),
	.parallelterminationcontrol_15(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ),
	.seriesterminationcontrol_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ),
	.seriesterminationcontrol_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ),
	.seriesterminationcontrol_2(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ),
	.seriesterminationcontrol_3(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ),
	.seriesterminationcontrol_4(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ),
	.seriesterminationcontrol_5(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ),
	.seriesterminationcontrol_6(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ),
	.seriesterminationcontrol_7(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ),
	.seriesterminationcontrol_8(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ),
	.seriesterminationcontrol_9(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ),
	.seriesterminationcontrol_10(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ),
	.seriesterminationcontrol_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ),
	.seriesterminationcontrol_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ),
	.seriesterminationcontrol_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ),
	.seriesterminationcontrol_14(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ),
	.seriesterminationcontrol_15(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ),
	.dqsin(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dataout_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ),
	.dataout_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ),
	.dataout_2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ),
	.dataout_3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ),
	.dataout_4(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ),
	.dataout_5(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ),
	.dataout_6(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ),
	.dataout_7(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ),
	.dataout_8(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ),
	.dataout_9(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ),
	.dataout_10(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ),
	.dataout_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ),
	.dataout_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ),
	.dataout_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ),
	.dataout_14(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ),
	.dataout_01(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ),
	.dataout_15(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ),
	.dataout_21(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ),
	.dataout_16(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ),
	.dataout_02(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ),
	.dataout_31(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ),
	.dataout_41(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ),
	.dataout_51(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ),
	.dataout_03(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ),
	.dataout_22(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ),
	.extra_output_pad_gen0delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.wire_pseudo_diffa_o_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.wire_pseudo_diffa_obar_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.wire_pseudo_diffa_oeout_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.wire_pseudo_diffa_oebout_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.pad_gen0delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.os(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.hps_io_emac1_inst_MDIO_0(\arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ),
	.hps_io_qspi_inst_IO0_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ),
	.hps_io_qspi_inst_IO1_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ),
	.hps_io_qspi_inst_IO2_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ),
	.hps_io_qspi_inst_IO3_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ),
	.hps_io_sdio_inst_CMD_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ),
	.hps_io_sdio_inst_D0_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ),
	.hps_io_sdio_inst_D1_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ),
	.hps_io_sdio_inst_D2_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ),
	.hps_io_sdio_inst_D3_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D0_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ),
	.hps_io_usb1_inst_D1_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ),
	.hps_io_usb1_inst_D2_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ),
	.hps_io_usb1_inst_D3_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D4_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ),
	.hps_io_usb1_inst_D5_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ),
	.hps_io_usb1_inst_D6_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ),
	.hps_io_usb1_inst_D7_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ),
	.hps_io_i2c0_inst_SDA_0(\arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o ),
	.hps_io_i2c0_inst_SCL_0(\arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o ),
	.hps_io_i2c1_inst_SDA_0(\arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o ),
	.hps_io_i2c1_inst_SCL_0(\arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o ),
	.hps_io_gpio_inst_GPIO09_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o ),
	.hps_io_gpio_inst_GPIO35_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~input_o ),
	.hps_io_gpio_inst_GPIO40_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o ),
	.hps_io_gpio_inst_GPIO41_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~input_o ),
	.hps_io_gpio_inst_GPIO48_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o ),
	.hps_io_gpio_inst_GPIO53_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~input_o ),
	.hps_io_gpio_inst_GPIO54_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~input_o ),
	.hps_io_gpio_inst_GPIO61_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o ),
	.hps_f2h_irq0_irq_0(\hps_f2h_irq0_irq[0]~input_o ),
	.hps_f2h_irq0_irq_1(\hps_f2h_irq0_irq[1]~input_o ),
	.hps_f2h_irq0_irq_2(\hps_f2h_irq0_irq[2]~input_o ),
	.hps_f2h_irq0_irq_3(\hps_f2h_irq0_irq[3]~input_o ),
	.hps_f2h_irq0_irq_4(\hps_f2h_irq0_irq[4]~input_o ),
	.hps_f2h_irq0_irq_5(\hps_f2h_irq0_irq[5]~input_o ),
	.hps_f2h_irq0_irq_6(\hps_f2h_irq0_irq[6]~input_o ),
	.hps_f2h_irq0_irq_7(\hps_f2h_irq0_irq[7]~input_o ),
	.hps_f2h_irq0_irq_8(\hps_f2h_irq0_irq[8]~input_o ),
	.hps_f2h_irq0_irq_9(\hps_f2h_irq0_irq[9]~input_o ),
	.hps_f2h_irq0_irq_10(\hps_f2h_irq0_irq[10]~input_o ),
	.hps_f2h_irq0_irq_11(\hps_f2h_irq0_irq[11]~input_o ),
	.hps_f2h_irq0_irq_12(\hps_f2h_irq0_irq[12]~input_o ),
	.hps_f2h_irq0_irq_13(\hps_f2h_irq0_irq[13]~input_o ),
	.hps_f2h_irq0_irq_14(\hps_f2h_irq0_irq[14]~input_o ),
	.hps_f2h_irq0_irq_15(\hps_f2h_irq0_irq[15]~input_o ),
	.hps_f2h_irq0_irq_16(\hps_f2h_irq0_irq[16]~input_o ),
	.hps_f2h_irq0_irq_17(\hps_f2h_irq0_irq[17]~input_o ),
	.hps_f2h_irq0_irq_18(\hps_f2h_irq0_irq[18]~input_o ),
	.hps_f2h_irq0_irq_19(\hps_f2h_irq0_irq[19]~input_o ),
	.hps_f2h_irq0_irq_20(\hps_f2h_irq0_irq[20]~input_o ),
	.hps_f2h_irq0_irq_21(\hps_f2h_irq0_irq[21]~input_o ),
	.hps_f2h_irq0_irq_22(\hps_f2h_irq0_irq[22]~input_o ),
	.hps_f2h_irq0_irq_23(\hps_f2h_irq0_irq[23]~input_o ),
	.hps_f2h_irq0_irq_24(\hps_f2h_irq0_irq[24]~input_o ),
	.hps_f2h_irq0_irq_25(\hps_f2h_irq0_irq[25]~input_o ),
	.hps_f2h_irq0_irq_26(\hps_f2h_irq0_irq[26]~input_o ),
	.hps_f2h_irq0_irq_27(\hps_f2h_irq0_irq[27]~input_o ),
	.hps_f2h_irq0_irq_28(\hps_f2h_irq0_irq[28]~input_o ),
	.hps_f2h_irq0_irq_29(\hps_f2h_irq0_irq[29]~input_o ),
	.hps_f2h_irq0_irq_30(\hps_f2h_irq0_irq[30]~input_o ),
	.hps_f2h_irq0_irq_31(\hps_f2h_irq0_irq[31]~input_o ),
	.hps_io_hps_io_emac1_inst_RXD0(\hps_io_hps_io_emac1_inst_RXD0~input_o ),
	.hps_io_hps_io_emac1_inst_RXD1(\hps_io_hps_io_emac1_inst_RXD1~input_o ),
	.hps_io_hps_io_emac1_inst_RXD2(\hps_io_hps_io_emac1_inst_RXD2~input_o ),
	.hps_io_hps_io_emac1_inst_RXD3(\hps_io_hps_io_emac1_inst_RXD3~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CLK(\hps_io_hps_io_emac1_inst_RX_CLK~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CTL(\hps_io_hps_io_emac1_inst_RX_CTL~input_o ),
	.hps_io_hps_io_spim1_inst_MISO(\hps_io_hps_io_spim1_inst_MISO~input_o ),
	.hps_io_hps_io_uart0_inst_RX(\hps_io_hps_io_uart0_inst_RX~input_o ),
	.hps_io_hps_io_usb1_inst_CLK(\hps_io_hps_io_usb1_inst_CLK~input_o ),
	.hps_io_hps_io_usb1_inst_DIR(\hps_io_hps_io_usb1_inst_DIR~input_o ),
	.hps_io_hps_io_usb1_inst_NXT(\hps_io_hps_io_usb1_inst_NXT~input_o ),
	.memory_oct_rzqin(\memory_oct_rzqin~input_o ));

Computer_System_Computer_System_mm_interconnect_0 mm_interconnect_0(
	.h2f_lw_ARVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARADDR_5(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[5] ),
	.h2f_lw_ARBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWADDR_5(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[5] ),
	.h2f_lw_AWBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.hold_waitrequest(\mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ),
	.WideOr0(\mm_interconnect_0|dma_2_control_port_slave_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|dma_2_control_port_slave_translator|wait_latency_counter[1]~q ),
	.WideOr01(\mm_interconnect_0|dma_1_control_port_slave_agent|WideOr0~0_combout ),
	.wait_latency_counter_11(\mm_interconnect_0|dma_1_control_port_slave_translator|wait_latency_counter[1]~q ),
	.cmd_sink_ready(\mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_rd_limiter|cmd_sink_ready~1_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.nonposted_cmd_accepted1(\mm_interconnect_0|arm_a9_hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ),
	.src_data_88(\mm_interconnect_0|rsp_mux|src_data[88]~combout ),
	.src_data_89(\mm_interconnect_0|rsp_mux|src_data[89]~combout ),
	.src_data_90(\mm_interconnect_0|rsp_mux|src_data[90]~combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux|src_data[91]~combout ),
	.src_data_92(\mm_interconnect_0|rsp_mux|src_data[92]~combout ),
	.src_data_93(\mm_interconnect_0|rsp_mux|src_data[93]~combout ),
	.src_data_94(\mm_interconnect_0|rsp_mux|src_data[94]~combout ),
	.src_data_95(\mm_interconnect_0|rsp_mux|src_data[95]~combout ),
	.src_data_96(\mm_interconnect_0|rsp_mux|src_data[96]~combout ),
	.src_data_97(\mm_interconnect_0|rsp_mux|src_data[97]~combout ),
	.src_data_98(\mm_interconnect_0|rsp_mux|src_data[98]~combout ),
	.src_data_99(\mm_interconnect_0|rsp_mux|src_data[99]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~2_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux_001|src_data[1]~5_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~8_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux_001|src_data[3]~11_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux_001|src_data[4]~14_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~17_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~20_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~23_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~26_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~29_combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~32_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[11]~35_combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~38_combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux_001|src_data[13]~41_combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~44_combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~47_combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~50_combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~53_combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~56_combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~59_combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux_001|src_data[20]~62_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[21]~65_combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~68_combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~71_combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~74_combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~77_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~80_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~83_combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~86_combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~89_combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~92_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[31]~95_combout ),
	.src_data_881(\mm_interconnect_0|rsp_mux_001|src_data[88]~combout ),
	.src_data_891(\mm_interconnect_0|rsp_mux_001|src_data[89]~combout ),
	.src_data_901(\mm_interconnect_0|rsp_mux_001|src_data[90]~combout ),
	.src_data_911(\mm_interconnect_0|rsp_mux_001|src_data[91]~combout ),
	.src_data_921(\mm_interconnect_0|rsp_mux_001|src_data[92]~combout ),
	.src_data_931(\mm_interconnect_0|rsp_mux_001|src_data[93]~combout ),
	.src_data_941(\mm_interconnect_0|rsp_mux_001|src_data[94]~combout ),
	.src_data_951(\mm_interconnect_0|rsp_mux_001|src_data[95]~combout ),
	.src_data_961(\mm_interconnect_0|rsp_mux_001|src_data[96]~combout ),
	.src_data_971(\mm_interconnect_0|rsp_mux_001|src_data[97]~combout ),
	.src_data_981(\mm_interconnect_0|rsp_mux_001|src_data[98]~combout ),
	.src_data_991(\mm_interconnect_0|rsp_mux_001|src_data[99]~combout ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.in_data_reg_2(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_59(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.mem(\mm_interconnect_0|dma_1_control_port_slave_agent_rsp_fifo|mem~0_combout ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_3(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.in_data_reg_210(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_591(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.mem1(\mm_interconnect_0|dma_2_control_port_slave_agent_rsp_fifo|mem~0_combout ),
	.int_nxt_addr_reg_dly_21(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_41(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_31(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_32(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_41(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_51(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_61(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_71(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_81(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_91(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_101(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_111(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_121(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_131(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_141(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_151(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_161(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_171(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_181(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_191(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_201(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_211(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_221(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_231(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_241(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_251(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_261(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_271(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_281(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_291(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_301(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_311(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.in_data_reg_0(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_1(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.dma_ctl_readdata_0(\dma_1|dma_ctl_readdata[0]~q ),
	.dma_ctl_readdata_01(\dma_2|dma_ctl_readdata[0]~q ),
	.dma_ctl_readdata_1(\dma_1|dma_ctl_readdata[1]~q ),
	.dma_ctl_readdata_11(\dma_2|dma_ctl_readdata[1]~q ),
	.dma_ctl_readdata_2(\dma_1|dma_ctl_readdata[2]~q ),
	.dma_ctl_readdata_21(\dma_2|dma_ctl_readdata[2]~q ),
	.dma_ctl_readdata_3(\dma_1|dma_ctl_readdata[3]~q ),
	.dma_ctl_readdata_31(\dma_2|dma_ctl_readdata[3]~q ),
	.dma_ctl_readdata_4(\dma_1|dma_ctl_readdata[4]~q ),
	.dma_ctl_readdata_41(\dma_2|dma_ctl_readdata[4]~q ),
	.dma_ctl_readdata_5(\dma_1|dma_ctl_readdata[5]~q ),
	.dma_ctl_readdata_51(\dma_2|dma_ctl_readdata[5]~q ),
	.dma_ctl_readdata_6(\dma_1|dma_ctl_readdata[6]~q ),
	.dma_ctl_readdata_61(\dma_2|dma_ctl_readdata[6]~q ),
	.dma_ctl_readdata_7(\dma_1|dma_ctl_readdata[7]~q ),
	.dma_ctl_readdata_71(\dma_2|dma_ctl_readdata[7]~q ),
	.dma_ctl_readdata_8(\dma_1|dma_ctl_readdata[8]~q ),
	.dma_ctl_readdata_81(\dma_2|dma_ctl_readdata[8]~q ),
	.dma_ctl_readdata_9(\dma_1|dma_ctl_readdata[9]~q ),
	.dma_ctl_readdata_91(\dma_2|dma_ctl_readdata[9]~q ),
	.dma_ctl_readdata_10(\dma_1|dma_ctl_readdata[10]~q ),
	.dma_ctl_readdata_101(\dma_2|dma_ctl_readdata[10]~q ),
	.dma_ctl_readdata_111(\dma_1|dma_ctl_readdata[11]~q ),
	.dma_ctl_readdata_112(\dma_2|dma_ctl_readdata[11]~q ),
	.dma_ctl_readdata_12(\dma_1|dma_ctl_readdata[12]~q ),
	.dma_ctl_readdata_121(\dma_2|dma_ctl_readdata[12]~q ),
	.dma_ctl_readdata_13(\dma_1|dma_ctl_readdata[13]~q ),
	.dma_ctl_readdata_131(\dma_2|dma_ctl_readdata[13]~q ),
	.dma_ctl_readdata_14(\dma_1|dma_ctl_readdata[14]~q ),
	.dma_ctl_readdata_141(\dma_2|dma_ctl_readdata[14]~q ),
	.dma_ctl_readdata_15(\dma_1|dma_ctl_readdata[15]~q ),
	.dma_ctl_readdata_151(\dma_2|dma_ctl_readdata[15]~q ),
	.dma_ctl_readdata_16(\dma_1|dma_ctl_readdata[16]~q ),
	.dma_ctl_readdata_161(\dma_2|dma_ctl_readdata[16]~q ),
	.dma_ctl_readdata_17(\dma_1|dma_ctl_readdata[17]~q ),
	.dma_ctl_readdata_171(\dma_2|dma_ctl_readdata[17]~q ),
	.dma_ctl_readdata_18(\dma_1|dma_ctl_readdata[18]~q ),
	.dma_ctl_readdata_181(\dma_2|dma_ctl_readdata[18]~q ),
	.dma_ctl_readdata_19(\dma_1|dma_ctl_readdata[19]~q ),
	.dma_ctl_readdata_191(\dma_2|dma_ctl_readdata[19]~q ),
	.dma_ctl_readdata_20(\dma_1|dma_ctl_readdata[20]~q ),
	.dma_ctl_readdata_201(\dma_2|dma_ctl_readdata[20]~q ),
	.dma_ctl_readdata_211(\dma_1|dma_ctl_readdata[21]~q ),
	.dma_ctl_readdata_212(\dma_2|dma_ctl_readdata[21]~q ),
	.dma_ctl_readdata_22(\dma_1|dma_ctl_readdata[22]~q ),
	.dma_ctl_readdata_221(\dma_2|dma_ctl_readdata[22]~q ),
	.dma_ctl_readdata_23(\dma_1|dma_ctl_readdata[23]~q ),
	.dma_ctl_readdata_231(\dma_2|dma_ctl_readdata[23]~q ),
	.dma_ctl_readdata_24(\dma_1|dma_ctl_readdata[24]~q ),
	.dma_ctl_readdata_241(\dma_2|dma_ctl_readdata[24]~q ),
	.dma_ctl_readdata_25(\dma_1|dma_ctl_readdata[25]~q ),
	.dma_ctl_readdata_251(\dma_2|dma_ctl_readdata[25]~q ),
	.dma_ctl_readdata_26(\dma_1|dma_ctl_readdata[26]~q ),
	.dma_ctl_readdata_261(\dma_2|dma_ctl_readdata[26]~q ),
	.dma_ctl_readdata_27(\dma_1|dma_ctl_readdata[27]~q ),
	.dma_ctl_readdata_271(\dma_2|dma_ctl_readdata[27]~q ),
	.dma_ctl_readdata_28(\dma_1|dma_ctl_readdata[28]~q ),
	.dma_ctl_readdata_281(\dma_2|dma_ctl_readdata[28]~q ),
	.dma_ctl_readdata_29(\dma_1|dma_ctl_readdata[29]~q ),
	.dma_ctl_readdata_291(\dma_2|dma_ctl_readdata[29]~q ),
	.dma_ctl_readdata_30(\dma_1|dma_ctl_readdata[30]~q ),
	.dma_ctl_readdata_301(\dma_2|dma_ctl_readdata[30]~q ),
	.dma_ctl_readdata_311(\dma_1|dma_ctl_readdata[31]~q ),
	.dma_ctl_readdata_312(\dma_2|dma_ctl_readdata[31]~q ),
	.in_data_reg_01(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_110(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ));

Computer_System_Computer_System_dma_2 dma_2(
	.f2h_AWREADY_0(\arm_a9_hps|fpga_interfaces|f2h_AWREADY[0] ),
	.f2h_WREADY_0(\arm_a9_hps|fpga_interfaces|f2h_WREADY[0] ),
	.ram_block1a32(\onchip_sram|the_altsyncram|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a0(\onchip_sram|the_altsyncram|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a33(\onchip_sram|the_altsyncram|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a1(\onchip_sram|the_altsyncram|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a34(\onchip_sram|the_altsyncram|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a2(\onchip_sram|the_altsyncram|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a35(\onchip_sram|the_altsyncram|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a3(\onchip_sram|the_altsyncram|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a36(\onchip_sram|the_altsyncram|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a4(\onchip_sram|the_altsyncram|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a37(\onchip_sram|the_altsyncram|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a5(\onchip_sram|the_altsyncram|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a38(\onchip_sram|the_altsyncram|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a6(\onchip_sram|the_altsyncram|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a39(\onchip_sram|the_altsyncram|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a7(\onchip_sram|the_altsyncram|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a40(\onchip_sram|the_altsyncram|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a8(\onchip_sram|the_altsyncram|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a41(\onchip_sram|the_altsyncram|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a9(\onchip_sram|the_altsyncram|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a42(\onchip_sram|the_altsyncram|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a10(\onchip_sram|the_altsyncram|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a43(\onchip_sram|the_altsyncram|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a11(\onchip_sram|the_altsyncram|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a44(\onchip_sram|the_altsyncram|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a12(\onchip_sram|the_altsyncram|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a45(\onchip_sram|the_altsyncram|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a13(\onchip_sram|the_altsyncram|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a46(\onchip_sram|the_altsyncram|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a14(\onchip_sram|the_altsyncram|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a47(\onchip_sram|the_altsyncram|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a15(\onchip_sram|the_altsyncram|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a56(\onchip_sram|the_altsyncram|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a24(\onchip_sram|the_altsyncram|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a57(\onchip_sram|the_altsyncram|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a25(\onchip_sram|the_altsyncram|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a58(\onchip_sram|the_altsyncram|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a26(\onchip_sram|the_altsyncram|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a59(\onchip_sram|the_altsyncram|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a27(\onchip_sram|the_altsyncram|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a60(\onchip_sram|the_altsyncram|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a28(\onchip_sram|the_altsyncram|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a61(\onchip_sram|the_altsyncram|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a29(\onchip_sram|the_altsyncram|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a62(\onchip_sram|the_altsyncram|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a30(\onchip_sram|the_altsyncram|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a63(\onchip_sram|the_altsyncram|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a31(\onchip_sram|the_altsyncram|auto_generated|ram_block1a31~portadataout ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.writeaddress_2(\dma_2|writeaddress[2]~q ),
	.writeaddress_3(\dma_2|writeaddress[3]~q ),
	.writeaddress_4(\dma_2|writeaddress[4]~q ),
	.writeaddress_5(\dma_2|writeaddress[5]~q ),
	.writeaddress_6(\dma_2|writeaddress[6]~q ),
	.writeaddress_7(\dma_2|writeaddress[7]~q ),
	.writeaddress_8(\dma_2|writeaddress[8]~q ),
	.writeaddress_9(\dma_2|writeaddress[9]~q ),
	.writeaddress_10(\dma_2|writeaddress[10]~q ),
	.writeaddress_11(\dma_2|writeaddress[11]~q ),
	.writeaddress_12(\dma_2|writeaddress[12]~q ),
	.writeaddress_13(\dma_2|writeaddress[13]~q ),
	.writeaddress_14(\dma_2|writeaddress[14]~q ),
	.writeaddress_15(\dma_2|writeaddress[15]~q ),
	.writeaddress_16(\dma_2|writeaddress[16]~q ),
	.writeaddress_17(\dma_2|writeaddress[17]~q ),
	.writeaddress_18(\dma_2|writeaddress[18]~q ),
	.writeaddress_19(\dma_2|writeaddress[19]~q ),
	.writeaddress_20(\dma_2|writeaddress[20]~q ),
	.writeaddress_21(\dma_2|writeaddress[21]~q ),
	.writeaddress_22(\dma_2|writeaddress[22]~q ),
	.writeaddress_23(\dma_2|writeaddress[23]~q ),
	.writeaddress_24(\dma_2|writeaddress[24]~q ),
	.writeaddress_25(\dma_2|writeaddress[25]~q ),
	.writeaddress_26(\dma_2|writeaddress[26]~q ),
	.writeaddress_27(\dma_2|writeaddress[27]~q ),
	.writeaddress_28(\dma_2|writeaddress[28]~q ),
	.writeaddress_29(\dma_2|writeaddress[29]~q ),
	.writeaddress_30(\dma_2|writeaddress[30]~q ),
	.writeaddress_31(\dma_2|writeaddress[31]~q ),
	.q_b_0(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[0] ),
	.q_b_1(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[1] ),
	.q_b_2(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[2] ),
	.q_b_3(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[3] ),
	.q_b_4(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[4] ),
	.q_b_5(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[5] ),
	.q_b_6(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[6] ),
	.q_b_7(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[7] ),
	.q_b_8(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[8] ),
	.q_b_9(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[9] ),
	.q_b_10(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[10] ),
	.q_b_11(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[11] ),
	.q_b_12(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[12] ),
	.q_b_13(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[13] ),
	.q_b_14(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[14] ),
	.q_b_15(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[15] ),
	.q_b_16(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[16] ),
	.q_b_17(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[17] ),
	.q_b_18(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[18] ),
	.q_b_19(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[19] ),
	.q_b_20(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[20] ),
	.q_b_21(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[21] ),
	.q_b_22(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[22] ),
	.q_b_23(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[23] ),
	.q_b_24(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[24] ),
	.q_b_25(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[25] ),
	.q_b_26(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[26] ),
	.q_b_27(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[27] ),
	.q_b_28(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[28] ),
	.q_b_29(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[29] ),
	.q_b_30(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[30] ),
	.q_b_31(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[31] ),
	.writeaddress_1(\dma_2|writeaddress[1]~q ),
	.writeaddress_0(\dma_2|writeaddress[0]~q ),
	.readaddress_15(\dma_2|readaddress[15]~q ),
	.readaddress_2(\dma_2|readaddress[2]~q ),
	.readaddress_3(\dma_2|readaddress[3]~q ),
	.readaddress_4(\dma_2|readaddress[4]~q ),
	.readaddress_5(\dma_2|readaddress[5]~q ),
	.readaddress_6(\dma_2|readaddress[6]~q ),
	.readaddress_7(\dma_2|readaddress[7]~q ),
	.readaddress_8(\dma_2|readaddress[8]~q ),
	.readaddress_9(\dma_2|readaddress[9]~q ),
	.readaddress_10(\dma_2|readaddress[10]~q ),
	.readaddress_11(\dma_2|readaddress[11]~q ),
	.readaddress_12(\dma_2|readaddress[12]~q ),
	.readaddress_13(\dma_2|readaddress[13]~q ),
	.readaddress_14(\dma_2|readaddress[14]~q ),
	.hold_waitrequest(\mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ),
	.address_taken(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|address_taken~q ),
	.mem_used_7(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[7]~q ),
	.fifo_empty(\dma_2|the_Computer_System_dma_2_fifo_module|fifo_empty~q ),
	.src_valid(\mm_interconnect_1|cmd_mux|src_valid~0_combout ),
	.data_taken(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|data_taken~q ),
	.last_write_collision(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_collision~q ),
	.last_write_data_0(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[0]~q ),
	.control_2(\dma_2|control[2]~q ),
	.control_0(\dma_2|control[0]~q ),
	.last_write_data_1(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[1]~q ),
	.last_write_data_2(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[2]~q ),
	.last_write_data_3(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[3]~q ),
	.last_write_data_4(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[4]~q ),
	.last_write_data_5(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[5]~q ),
	.last_write_data_6(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[6]~q ),
	.last_write_data_7(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[7]~q ),
	.write_writedata(\dma_2|write_writedata~0_combout ),
	.last_write_data_8(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[8]~q ),
	.write_writedata1(\dma_2|write_writedata~1_combout ),
	.last_write_data_9(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[9]~q ),
	.write_writedata2(\dma_2|write_writedata~2_combout ),
	.last_write_data_10(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[10]~q ),
	.write_writedata3(\dma_2|write_writedata~3_combout ),
	.last_write_data_11(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[11]~q ),
	.write_writedata4(\dma_2|write_writedata~4_combout ),
	.last_write_data_12(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[12]~q ),
	.write_writedata5(\dma_2|write_writedata~5_combout ),
	.last_write_data_13(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[13]~q ),
	.write_writedata6(\dma_2|write_writedata~6_combout ),
	.last_write_data_14(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[14]~q ),
	.write_writedata7(\dma_2|write_writedata~7_combout ),
	.last_write_data_15(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[15]~q ),
	.last_write_data_16(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[16]~q ),
	.last_write_data_17(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[17]~q ),
	.last_write_data_18(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[18]~q ),
	.last_write_data_19(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[19]~q ),
	.last_write_data_20(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[20]~q ),
	.last_write_data_21(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[21]~q ),
	.last_write_data_22(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[22]~q ),
	.last_write_data_23(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[23]~q ),
	.last_write_data_24(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[24]~q ),
	.last_write_data_25(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[25]~q ),
	.last_write_data_26(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[26]~q ),
	.last_write_data_27(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[27]~q ),
	.last_write_data_28(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[28]~q ),
	.last_write_data_29(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[29]~q ),
	.last_write_data_30(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[30]~q ),
	.last_write_data_31(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[31]~q ),
	.WideOr0(\mm_interconnect_0|dma_2_control_port_slave_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|dma_2_control_port_slave_translator|wait_latency_counter[1]~q ),
	.saved_grant_0(\mm_interconnect_2|cmd_mux|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_2|onchip_sram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.system_reset_n(\rst_controller|r_sync_rst~q ),
	.fifo_read(\dma_2|the_Computer_System_dma_2_mem_write|fifo_read~0_combout ),
	.write_cp_ready(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|write_cp_ready~0_combout ),
	.src0_valid(\mm_interconnect_2|rsp_demux|src0_valid~combout ),
	.in_data_reg_2(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_59(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.mem(\mm_interconnect_0|dma_2_control_port_slave_agent_rsp_fifo|mem~0_combout ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_3(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.address_reg_a_0(\onchip_sram|the_altsyncram|auto_generated|address_reg_a[0]~q ),
	.l1_w16_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w16_n0_mux_dataout~0_combout ),
	.in_data_reg_0(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.l1_w17_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w17_n0_mux_dataout~0_combout ),
	.l1_w18_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w18_n0_mux_dataout~0_combout ),
	.l1_w19_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w19_n0_mux_dataout~0_combout ),
	.l1_w20_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w20_n0_mux_dataout~0_combout ),
	.l1_w21_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w21_n0_mux_dataout~0_combout ),
	.l1_w22_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w22_n0_mux_dataout~0_combout ),
	.l1_w23_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w23_n0_mux_dataout~0_combout ),
	.l1_w8_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w8_n0_mux_dataout~0_combout ),
	.l1_w9_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w9_n0_mux_dataout~0_combout ),
	.l1_w10_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w10_n0_mux_dataout~0_combout ),
	.l1_w11_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w11_n0_mux_dataout~0_combout ),
	.l1_w12_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w12_n0_mux_dataout~0_combout ),
	.l1_w13_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w13_n0_mux_dataout~0_combout ),
	.l1_w14_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w14_n0_mux_dataout~0_combout ),
	.l1_w15_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w15_n0_mux_dataout~0_combout ),
	.l1_w24_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w24_n0_mux_dataout~0_combout ),
	.l1_w25_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w25_n0_mux_dataout~0_combout ),
	.l1_w26_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w26_n0_mux_dataout~0_combout ),
	.l1_w27_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w27_n0_mux_dataout~0_combout ),
	.l1_w28_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w28_n0_mux_dataout~0_combout ),
	.l1_w29_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w29_n0_mux_dataout~0_combout ),
	.l1_w30_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w30_n0_mux_dataout~0_combout ),
	.l1_w31_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w31_n0_mux_dataout~0_combout ),
	.in_data_reg_1(\mm_interconnect_0|dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.dma_ctl_readdata_0(\dma_2|dma_ctl_readdata[0]~q ),
	.dma_ctl_readdata_1(\dma_2|dma_ctl_readdata[1]~q ),
	.dma_ctl_readdata_2(\dma_2|dma_ctl_readdata[2]~q ),
	.dma_ctl_readdata_3(\dma_2|dma_ctl_readdata[3]~q ),
	.dma_ctl_readdata_4(\dma_2|dma_ctl_readdata[4]~q ),
	.dma_ctl_readdata_5(\dma_2|dma_ctl_readdata[5]~q ),
	.dma_ctl_readdata_6(\dma_2|dma_ctl_readdata[6]~q ),
	.dma_ctl_readdata_7(\dma_2|dma_ctl_readdata[7]~q ),
	.dma_ctl_readdata_8(\dma_2|dma_ctl_readdata[8]~q ),
	.dma_ctl_readdata_9(\dma_2|dma_ctl_readdata[9]~q ),
	.dma_ctl_readdata_10(\dma_2|dma_ctl_readdata[10]~q ),
	.dma_ctl_readdata_11(\dma_2|dma_ctl_readdata[11]~q ),
	.dma_ctl_readdata_12(\dma_2|dma_ctl_readdata[12]~q ),
	.dma_ctl_readdata_13(\dma_2|dma_ctl_readdata[13]~q ),
	.dma_ctl_readdata_14(\dma_2|dma_ctl_readdata[14]~q ),
	.dma_ctl_readdata_15(\dma_2|dma_ctl_readdata[15]~q ),
	.dma_ctl_readdata_16(\dma_2|dma_ctl_readdata[16]~q ),
	.dma_ctl_readdata_17(\dma_2|dma_ctl_readdata[17]~q ),
	.dma_ctl_readdata_18(\dma_2|dma_ctl_readdata[18]~q ),
	.dma_ctl_readdata_19(\dma_2|dma_ctl_readdata[19]~q ),
	.dma_ctl_readdata_20(\dma_2|dma_ctl_readdata[20]~q ),
	.dma_ctl_readdata_21(\dma_2|dma_ctl_readdata[21]~q ),
	.dma_ctl_readdata_22(\dma_2|dma_ctl_readdata[22]~q ),
	.dma_ctl_readdata_23(\dma_2|dma_ctl_readdata[23]~q ),
	.dma_ctl_readdata_24(\dma_2|dma_ctl_readdata[24]~q ),
	.dma_ctl_readdata_25(\dma_2|dma_ctl_readdata[25]~q ),
	.dma_ctl_readdata_26(\dma_2|dma_ctl_readdata[26]~q ),
	.dma_ctl_readdata_27(\dma_2|dma_ctl_readdata[27]~q ),
	.dma_ctl_readdata_28(\dma_2|dma_ctl_readdata[28]~q ),
	.dma_ctl_readdata_29(\dma_2|dma_ctl_readdata[29]~q ),
	.dma_ctl_readdata_30(\dma_2|dma_ctl_readdata[30]~q ),
	.dma_ctl_readdata_31(\dma_2|dma_ctl_readdata[31]~q ),
	.read_select(\dma_2|the_Computer_System_dma_2_mem_read|read_select~q ),
	.read_latency_shift_reg(\mm_interconnect_2|onchip_sram_s1_translator|read_latency_shift_reg~0_combout ));

Computer_System_Computer_System_Onchip_SRAM onchip_sram(
	.ram_block1a32(\onchip_sram|the_altsyncram|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a0(\onchip_sram|the_altsyncram|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a33(\onchip_sram|the_altsyncram|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a1(\onchip_sram|the_altsyncram|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a34(\onchip_sram|the_altsyncram|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a2(\onchip_sram|the_altsyncram|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a35(\onchip_sram|the_altsyncram|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a3(\onchip_sram|the_altsyncram|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a36(\onchip_sram|the_altsyncram|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a4(\onchip_sram|the_altsyncram|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a37(\onchip_sram|the_altsyncram|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a5(\onchip_sram|the_altsyncram|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a38(\onchip_sram|the_altsyncram|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a6(\onchip_sram|the_altsyncram|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a39(\onchip_sram|the_altsyncram|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a7(\onchip_sram|the_altsyncram|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a40(\onchip_sram|the_altsyncram|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a8(\onchip_sram|the_altsyncram|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a41(\onchip_sram|the_altsyncram|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a9(\onchip_sram|the_altsyncram|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a42(\onchip_sram|the_altsyncram|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a10(\onchip_sram|the_altsyncram|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a43(\onchip_sram|the_altsyncram|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a11(\onchip_sram|the_altsyncram|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a44(\onchip_sram|the_altsyncram|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a12(\onchip_sram|the_altsyncram|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a45(\onchip_sram|the_altsyncram|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a13(\onchip_sram|the_altsyncram|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a46(\onchip_sram|the_altsyncram|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a14(\onchip_sram|the_altsyncram|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a47(\onchip_sram|the_altsyncram|auto_generated|ram_block1a47~portadataout ),
	.ram_block1a15(\onchip_sram|the_altsyncram|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a56(\onchip_sram|the_altsyncram|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a24(\onchip_sram|the_altsyncram|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a57(\onchip_sram|the_altsyncram|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a25(\onchip_sram|the_altsyncram|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a58(\onchip_sram|the_altsyncram|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a26(\onchip_sram|the_altsyncram|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a59(\onchip_sram|the_altsyncram|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a27(\onchip_sram|the_altsyncram|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a60(\onchip_sram|the_altsyncram|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a28(\onchip_sram|the_altsyncram|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a61(\onchip_sram|the_altsyncram|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a29(\onchip_sram|the_altsyncram|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a62(\onchip_sram|the_altsyncram|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a30(\onchip_sram|the_altsyncram|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a63(\onchip_sram|the_altsyncram|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a31(\onchip_sram|the_altsyncram|auto_generated|ram_block1a31~portadataout ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.readaddress_15(\dma_2|readaddress[15]~q ),
	.writeaddress_15(\dma_1|writeaddress[15]~q ),
	.l1_w0_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w0_n0_mux_dataout~0_combout ),
	.l1_w1_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w1_n0_mux_dataout~0_combout ),
	.l1_w2_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w2_n0_mux_dataout~0_combout ),
	.l1_w3_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w3_n0_mux_dataout~0_combout ),
	.l1_w4_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w4_n0_mux_dataout~0_combout ),
	.l1_w5_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w5_n0_mux_dataout~0_combout ),
	.l1_w6_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w6_n0_mux_dataout~0_combout ),
	.l1_w7_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w7_n0_mux_dataout~0_combout ),
	.l1_w8_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w8_n0_mux_dataout~0_combout ),
	.l1_w9_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w9_n0_mux_dataout~0_combout ),
	.l1_w10_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w10_n0_mux_dataout~0_combout ),
	.l1_w11_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w11_n0_mux_dataout~0_combout ),
	.l1_w12_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w12_n0_mux_dataout~0_combout ),
	.l1_w13_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w13_n0_mux_dataout~0_combout ),
	.l1_w14_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w14_n0_mux_dataout~0_combout ),
	.l1_w15_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w15_n0_mux_dataout~0_combout ),
	.l1_w16_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w16_n0_mux_dataout~0_combout ),
	.l1_w17_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w17_n0_mux_dataout~0_combout ),
	.l1_w18_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w18_n0_mux_dataout~0_combout ),
	.l1_w19_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w19_n0_mux_dataout~0_combout ),
	.l1_w20_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w20_n0_mux_dataout~0_combout ),
	.l1_w21_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w21_n0_mux_dataout~0_combout ),
	.l1_w22_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w22_n0_mux_dataout~0_combout ),
	.l1_w23_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w23_n0_mux_dataout~0_combout ),
	.l1_w24_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w24_n0_mux_dataout~0_combout ),
	.l1_w25_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w25_n0_mux_dataout~0_combout ),
	.l1_w26_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w26_n0_mux_dataout~0_combout ),
	.l1_w27_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w27_n0_mux_dataout~0_combout ),
	.l1_w28_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w28_n0_mux_dataout~0_combout ),
	.l1_w29_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w29_n0_mux_dataout~0_combout ),
	.l1_w30_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w30_n0_mux_dataout~0_combout ),
	.l1_w31_n0_mux_dataout(\onchip_sram|the_altsyncram|auto_generated|mux5|l1_w31_n0_mux_dataout~0_combout ),
	.hold_waitrequest(\mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ),
	.saved_grant_0(\mm_interconnect_2|cmd_mux|saved_grant[0]~q ),
	.saved_grant_1(\mm_interconnect_2|cmd_mux|saved_grant[1]~q ),
	.mem_used_1(\mm_interconnect_2|onchip_sram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.fifo_empty(\dma_1|the_Computer_System_dma_1_fifo_module|fifo_empty~q ),
	.wren(\onchip_sram|wren~0_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_2|cmd_mux|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_2|cmd_mux|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_2|cmd_mux|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_2|cmd_mux|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_2|cmd_mux|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_2|cmd_mux|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_2|cmd_mux|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_2|cmd_mux|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_2|cmd_mux|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_2|cmd_mux|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_2|cmd_mux|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_2|cmd_mux|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_2|cmd_mux|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_2|cmd_mux|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_2|cmd_mux|src_data[32]~0_combout ),
	.src_payload1(\mm_interconnect_2|cmd_mux|src_payload~2_combout ),
	.src_payload2(\mm_interconnect_2|cmd_mux|src_payload~3_combout ),
	.src_payload3(\mm_interconnect_2|cmd_mux|src_payload~4_combout ),
	.src_payload4(\mm_interconnect_2|cmd_mux|src_payload~5_combout ),
	.src_payload5(\mm_interconnect_2|cmd_mux|src_payload~6_combout ),
	.src_payload6(\mm_interconnect_2|cmd_mux|src_payload~7_combout ),
	.src_payload7(\mm_interconnect_2|cmd_mux|src_payload~8_combout ),
	.src_payload8(\mm_interconnect_2|cmd_mux|src_payload~9_combout ),
	.src_data_33(\mm_interconnect_2|cmd_mux|src_data[33]~1_combout ),
	.src_payload9(\mm_interconnect_2|cmd_mux|src_payload~10_combout ),
	.src_payload10(\mm_interconnect_2|cmd_mux|src_payload~11_combout ),
	.src_payload11(\mm_interconnect_2|cmd_mux|src_payload~12_combout ),
	.src_payload12(\mm_interconnect_2|cmd_mux|src_payload~13_combout ),
	.src_payload13(\mm_interconnect_2|cmd_mux|src_payload~14_combout ),
	.src_payload14(\mm_interconnect_2|cmd_mux|src_payload~15_combout ),
	.src_payload15(\mm_interconnect_2|cmd_mux|src_payload~16_combout ),
	.src_payload16(\mm_interconnect_2|cmd_mux|src_payload~17_combout ),
	.src_data_34(\mm_interconnect_2|cmd_mux|src_data[34]~2_combout ),
	.src_payload17(\mm_interconnect_2|cmd_mux|src_payload~18_combout ),
	.src_payload18(\mm_interconnect_2|cmd_mux|src_payload~19_combout ),
	.src_payload19(\mm_interconnect_2|cmd_mux|src_payload~20_combout ),
	.src_payload20(\mm_interconnect_2|cmd_mux|src_payload~21_combout ),
	.src_payload21(\mm_interconnect_2|cmd_mux|src_payload~22_combout ),
	.src_payload22(\mm_interconnect_2|cmd_mux|src_payload~23_combout ),
	.src_payload23(\mm_interconnect_2|cmd_mux|src_payload~24_combout ),
	.src_payload24(\mm_interconnect_2|cmd_mux|src_payload~25_combout ),
	.src_data_35(\mm_interconnect_2|cmd_mux|src_data[35]~3_combout ),
	.src_payload25(\mm_interconnect_2|cmd_mux|src_payload~26_combout ),
	.src_payload26(\mm_interconnect_2|cmd_mux|src_payload~27_combout ),
	.src_payload27(\mm_interconnect_2|cmd_mux|src_payload~28_combout ),
	.src_payload28(\mm_interconnect_2|cmd_mux|src_payload~29_combout ),
	.src_payload29(\mm_interconnect_2|cmd_mux|src_payload~30_combout ),
	.src_payload30(\mm_interconnect_2|cmd_mux|src_payload~31_combout ),
	.src_payload31(\mm_interconnect_2|cmd_mux|src_payload~32_combout ),
	.address_reg_a_0(\onchip_sram|the_altsyncram|auto_generated|address_reg_a[0]~q ),
	.l1_w16_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w16_n0_mux_dataout~0_combout ),
	.l1_w17_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w17_n0_mux_dataout~0_combout ),
	.l1_w18_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w18_n0_mux_dataout~0_combout ),
	.l1_w19_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w19_n0_mux_dataout~0_combout ),
	.l1_w20_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w20_n0_mux_dataout~0_combout ),
	.l1_w21_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w21_n0_mux_dataout~0_combout ),
	.l1_w22_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w22_n0_mux_dataout~0_combout ),
	.l1_w23_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w23_n0_mux_dataout~0_combout ),
	.l1_w8_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w8_n0_mux_dataout~0_combout ),
	.l1_w9_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w9_n0_mux_dataout~0_combout ),
	.l1_w10_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w10_n0_mux_dataout~0_combout ),
	.l1_w11_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w11_n0_mux_dataout~0_combout ),
	.l1_w12_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w12_n0_mux_dataout~0_combout ),
	.l1_w13_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w13_n0_mux_dataout~0_combout ),
	.l1_w14_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w14_n0_mux_dataout~0_combout ),
	.l1_w15_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w15_n0_mux_dataout~0_combout ),
	.l1_w24_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w24_n0_mux_dataout~0_combout ),
	.l1_w25_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w25_n0_mux_dataout~0_combout ),
	.l1_w26_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w26_n0_mux_dataout~0_combout ),
	.l1_w27_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w27_n0_mux_dataout~0_combout ),
	.l1_w28_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w28_n0_mux_dataout~0_combout ),
	.l1_w29_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w29_n0_mux_dataout~0_combout ),
	.l1_w30_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w30_n0_mux_dataout~0_combout ),
	.l1_w31_n0_mux_dataout1(\onchip_sram|the_altsyncram|auto_generated|mux4|l1_w31_n0_mux_dataout~0_combout ),
	.src_data_51(\mm_interconnect_2|cmd_mux|src_data[51]~combout ),
	.onchip_sram_s2_address_13(\onchip_sram_s2_address[13]~input_o ),
	.onchip_sram_s2_chipselect(\onchip_sram_s2_chipselect~input_o ),
	.onchip_sram_s2_write(\onchip_sram_s2_write~input_o ),
	.onchip_sram_clk2_clk(\onchip_sram_clk2_clk~input_o ),
	.onchip_sram_reset2_reset_req(\onchip_sram_reset2_reset_req~input_o ),
	.onchip_sram_s2_clken(\onchip_sram_s2_clken~input_o ),
	.onchip_sram_s2_writedata_0(\onchip_sram_s2_writedata[0]~input_o ),
	.onchip_sram_s2_address_0(\onchip_sram_s2_address[0]~input_o ),
	.onchip_sram_s2_address_1(\onchip_sram_s2_address[1]~input_o ),
	.onchip_sram_s2_address_2(\onchip_sram_s2_address[2]~input_o ),
	.onchip_sram_s2_address_3(\onchip_sram_s2_address[3]~input_o ),
	.onchip_sram_s2_address_4(\onchip_sram_s2_address[4]~input_o ),
	.onchip_sram_s2_address_5(\onchip_sram_s2_address[5]~input_o ),
	.onchip_sram_s2_address_6(\onchip_sram_s2_address[6]~input_o ),
	.onchip_sram_s2_address_7(\onchip_sram_s2_address[7]~input_o ),
	.onchip_sram_s2_address_8(\onchip_sram_s2_address[8]~input_o ),
	.onchip_sram_s2_address_9(\onchip_sram_s2_address[9]~input_o ),
	.onchip_sram_s2_address_10(\onchip_sram_s2_address[10]~input_o ),
	.onchip_sram_s2_address_11(\onchip_sram_s2_address[11]~input_o ),
	.onchip_sram_s2_address_12(\onchip_sram_s2_address[12]~input_o ),
	.onchip_sram_s2_byteenable_0(\onchip_sram_s2_byteenable[0]~input_o ),
	.onchip_sram_s2_writedata_1(\onchip_sram_s2_writedata[1]~input_o ),
	.onchip_sram_s2_writedata_2(\onchip_sram_s2_writedata[2]~input_o ),
	.onchip_sram_s2_writedata_3(\onchip_sram_s2_writedata[3]~input_o ),
	.onchip_sram_s2_writedata_4(\onchip_sram_s2_writedata[4]~input_o ),
	.onchip_sram_s2_writedata_5(\onchip_sram_s2_writedata[5]~input_o ),
	.onchip_sram_s2_writedata_6(\onchip_sram_s2_writedata[6]~input_o ),
	.onchip_sram_s2_writedata_7(\onchip_sram_s2_writedata[7]~input_o ),
	.onchip_sram_s2_writedata_8(\onchip_sram_s2_writedata[8]~input_o ),
	.onchip_sram_s2_byteenable_1(\onchip_sram_s2_byteenable[1]~input_o ),
	.onchip_sram_s2_writedata_9(\onchip_sram_s2_writedata[9]~input_o ),
	.onchip_sram_s2_writedata_10(\onchip_sram_s2_writedata[10]~input_o ),
	.onchip_sram_s2_writedata_11(\onchip_sram_s2_writedata[11]~input_o ),
	.onchip_sram_s2_writedata_12(\onchip_sram_s2_writedata[12]~input_o ),
	.onchip_sram_s2_writedata_13(\onchip_sram_s2_writedata[13]~input_o ),
	.onchip_sram_s2_writedata_14(\onchip_sram_s2_writedata[14]~input_o ),
	.onchip_sram_s2_writedata_15(\onchip_sram_s2_writedata[15]~input_o ),
	.onchip_sram_s2_writedata_16(\onchip_sram_s2_writedata[16]~input_o ),
	.onchip_sram_s2_byteenable_2(\onchip_sram_s2_byteenable[2]~input_o ),
	.onchip_sram_s2_writedata_17(\onchip_sram_s2_writedata[17]~input_o ),
	.onchip_sram_s2_writedata_18(\onchip_sram_s2_writedata[18]~input_o ),
	.onchip_sram_s2_writedata_19(\onchip_sram_s2_writedata[19]~input_o ),
	.onchip_sram_s2_writedata_20(\onchip_sram_s2_writedata[20]~input_o ),
	.onchip_sram_s2_writedata_21(\onchip_sram_s2_writedata[21]~input_o ),
	.onchip_sram_s2_writedata_22(\onchip_sram_s2_writedata[22]~input_o ),
	.onchip_sram_s2_writedata_23(\onchip_sram_s2_writedata[23]~input_o ),
	.onchip_sram_s2_writedata_24(\onchip_sram_s2_writedata[24]~input_o ),
	.onchip_sram_s2_byteenable_3(\onchip_sram_s2_byteenable[3]~input_o ),
	.onchip_sram_s2_writedata_25(\onchip_sram_s2_writedata[25]~input_o ),
	.onchip_sram_s2_writedata_26(\onchip_sram_s2_writedata[26]~input_o ),
	.onchip_sram_s2_writedata_27(\onchip_sram_s2_writedata[27]~input_o ),
	.onchip_sram_s2_writedata_28(\onchip_sram_s2_writedata[28]~input_o ),
	.onchip_sram_s2_writedata_29(\onchip_sram_s2_writedata[29]~input_o ),
	.onchip_sram_s2_writedata_30(\onchip_sram_s2_writedata[30]~input_o ),
	.onchip_sram_s2_writedata_31(\onchip_sram_s2_writedata[31]~input_o ));

Computer_System_Computer_System_dma_1 dma_1(
	.f2h_ARREADY_0(\arm_a9_hps|fpga_interfaces|f2h_ARREADY[0] ),
	.f2h_RVALID_0(\arm_a9_hps|fpga_interfaces|f2h_RVALID[0] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.readaddress_2(\dma_1|readaddress[2]~q ),
	.readaddress_3(\dma_1|readaddress[3]~q ),
	.readaddress_4(\dma_1|readaddress[4]~q ),
	.readaddress_5(\dma_1|readaddress[5]~q ),
	.readaddress_6(\dma_1|readaddress[6]~q ),
	.readaddress_7(\dma_1|readaddress[7]~q ),
	.readaddress_8(\dma_1|readaddress[8]~q ),
	.readaddress_9(\dma_1|readaddress[9]~q ),
	.readaddress_10(\dma_1|readaddress[10]~q ),
	.readaddress_11(\dma_1|readaddress[11]~q ),
	.readaddress_12(\dma_1|readaddress[12]~q ),
	.readaddress_13(\dma_1|readaddress[13]~q ),
	.readaddress_14(\dma_1|readaddress[14]~q ),
	.readaddress_15(\dma_1|readaddress[15]~q ),
	.readaddress_16(\dma_1|readaddress[16]~q ),
	.readaddress_17(\dma_1|readaddress[17]~q ),
	.readaddress_18(\dma_1|readaddress[18]~q ),
	.readaddress_19(\dma_1|readaddress[19]~q ),
	.readaddress_20(\dma_1|readaddress[20]~q ),
	.readaddress_21(\dma_1|readaddress[21]~q ),
	.readaddress_22(\dma_1|readaddress[22]~q ),
	.readaddress_23(\dma_1|readaddress[23]~q ),
	.readaddress_24(\dma_1|readaddress[24]~q ),
	.readaddress_25(\dma_1|readaddress[25]~q ),
	.readaddress_26(\dma_1|readaddress[26]~q ),
	.readaddress_27(\dma_1|readaddress[27]~q ),
	.readaddress_28(\dma_1|readaddress[28]~q ),
	.readaddress_29(\dma_1|readaddress[29]~q ),
	.readaddress_30(\dma_1|readaddress[30]~q ),
	.readaddress_31(\dma_1|readaddress[31]~q ),
	.writeaddress_15(\dma_1|writeaddress[15]~q ),
	.q_b_0(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[0] ),
	.writeaddress_2(\dma_1|writeaddress[2]~q ),
	.writeaddress_3(\dma_1|writeaddress[3]~q ),
	.writeaddress_4(\dma_1|writeaddress[4]~q ),
	.writeaddress_5(\dma_1|writeaddress[5]~q ),
	.writeaddress_6(\dma_1|writeaddress[6]~q ),
	.writeaddress_7(\dma_1|writeaddress[7]~q ),
	.writeaddress_8(\dma_1|writeaddress[8]~q ),
	.writeaddress_9(\dma_1|writeaddress[9]~q ),
	.writeaddress_10(\dma_1|writeaddress[10]~q ),
	.writeaddress_11(\dma_1|writeaddress[11]~q ),
	.writeaddress_12(\dma_1|writeaddress[12]~q ),
	.writeaddress_13(\dma_1|writeaddress[13]~q ),
	.writeaddress_14(\dma_1|writeaddress[14]~q ),
	.writeaddress_1(\dma_1|writeaddress[1]~q ),
	.writeaddress_0(\dma_1|writeaddress[0]~q ),
	.q_b_1(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[1] ),
	.q_b_2(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[2] ),
	.q_b_3(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[3] ),
	.q_b_4(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[4] ),
	.q_b_5(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[5] ),
	.q_b_6(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[6] ),
	.q_b_7(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[7] ),
	.q_b_8(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[8] ),
	.q_b_9(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[9] ),
	.q_b_10(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[10] ),
	.q_b_11(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[11] ),
	.q_b_12(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[12] ),
	.q_b_13(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[13] ),
	.q_b_14(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[14] ),
	.q_b_15(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[15] ),
	.q_b_16(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[16] ),
	.q_b_17(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[17] ),
	.q_b_18(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[18] ),
	.q_b_19(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[19] ),
	.q_b_20(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[20] ),
	.q_b_21(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[21] ),
	.q_b_22(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[22] ),
	.q_b_23(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[23] ),
	.q_b_24(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[24] ),
	.q_b_25(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[25] ),
	.q_b_26(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[26] ),
	.q_b_27(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[27] ),
	.q_b_28(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[28] ),
	.q_b_29(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[29] ),
	.q_b_30(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[30] ),
	.q_b_31(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[31] ),
	.mem_used_7(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem_used[7]~q ),
	.saved_grant_0(\mm_interconnect_1|cmd_mux_001|saved_grant[0]~q ),
	.read_select(\dma_1|the_Computer_System_dma_1_mem_read|read_select~q ),
	.hold_waitrequest(\mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ),
	.write(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|write~0_combout ),
	.WideOr0(\mm_interconnect_0|dma_1_control_port_slave_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|dma_1_control_port_slave_translator|wait_latency_counter[1]~q ),
	.saved_grant_1(\mm_interconnect_2|cmd_mux|saved_grant[1]~q ),
	.mem_used_1(\mm_interconnect_2|onchip_sram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.fifo_empty(\dma_1|the_Computer_System_dma_1_fifo_module|fifo_empty~q ),
	.wren(\onchip_sram|wren~0_combout ),
	.last_write_collision(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_collision~q ),
	.last_write_data_0(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[0]~q ),
	.control_2(\dma_1|control[2]~q ),
	.control_0(\dma_1|control[0]~q ),
	.last_write_data_1(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[1]~q ),
	.last_write_data_2(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[2]~q ),
	.last_write_data_3(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[3]~q ),
	.last_write_data_4(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[4]~q ),
	.last_write_data_5(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[5]~q ),
	.last_write_data_6(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[6]~q ),
	.last_write_data_7(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[7]~q ),
	.write_writedata(\dma_1|write_writedata~0_combout ),
	.last_write_data_8(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[8]~q ),
	.write_writedata1(\dma_1|write_writedata~1_combout ),
	.last_write_data_9(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[9]~q ),
	.write_writedata2(\dma_1|write_writedata~2_combout ),
	.last_write_data_10(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[10]~q ),
	.write_writedata3(\dma_1|write_writedata~3_combout ),
	.last_write_data_11(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[11]~q ),
	.write_writedata4(\dma_1|write_writedata~4_combout ),
	.last_write_data_12(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[12]~q ),
	.write_writedata5(\dma_1|write_writedata~5_combout ),
	.last_write_data_13(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[13]~q ),
	.write_writedata6(\dma_1|write_writedata~6_combout ),
	.last_write_data_14(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[14]~q ),
	.write_writedata7(\dma_1|write_writedata~7_combout ),
	.last_write_data_15(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[15]~q ),
	.last_write_data_16(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[16]~q ),
	.last_write_data_17(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[17]~q ),
	.last_write_data_18(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[18]~q ),
	.last_write_data_19(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[19]~q ),
	.last_write_data_20(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[20]~q ),
	.last_write_data_21(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[21]~q ),
	.last_write_data_22(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[22]~q ),
	.last_write_data_23(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[23]~q ),
	.last_write_data_24(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[24]~q ),
	.last_write_data_25(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[25]~q ),
	.last_write_data_26(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[26]~q ),
	.last_write_data_27(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[27]~q ),
	.last_write_data_28(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[28]~q ),
	.last_write_data_29(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[29]~q ),
	.last_write_data_30(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[30]~q ),
	.last_write_data_31(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[31]~q ),
	.WideOr1(\mm_interconnect_1|cmd_mux_001|WideOr1~0_combout ),
	.system_reset_n(\rst_controller|r_sync_rst~q ),
	.inc_read(\dma_1|the_Computer_System_dma_1_mem_read|inc_read~combout ),
	.av_readdatavalid(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~0_combout ),
	.av_readdatavalid1(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~1_combout ),
	.av_readdatavalid2(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~2_combout ),
	.av_readdatavalid3(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~3_combout ),
	.in_data_reg_2(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_59(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.mem(\mm_interconnect_0|dma_1_control_port_slave_agent_rsp_fifo|mem~0_combout ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_3(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.dma_ctl_readdata_0(\dma_1|dma_ctl_readdata[0]~q ),
	.dma_ctl_readdata_1(\dma_1|dma_ctl_readdata[1]~q ),
	.dma_ctl_readdata_2(\dma_1|dma_ctl_readdata[2]~q ),
	.dma_ctl_readdata_3(\dma_1|dma_ctl_readdata[3]~q ),
	.dma_ctl_readdata_4(\dma_1|dma_ctl_readdata[4]~q ),
	.dma_ctl_readdata_5(\dma_1|dma_ctl_readdata[5]~q ),
	.dma_ctl_readdata_6(\dma_1|dma_ctl_readdata[6]~q ),
	.dma_ctl_readdata_7(\dma_1|dma_ctl_readdata[7]~q ),
	.dma_ctl_readdata_8(\dma_1|dma_ctl_readdata[8]~q ),
	.dma_ctl_readdata_9(\dma_1|dma_ctl_readdata[9]~q ),
	.dma_ctl_readdata_10(\dma_1|dma_ctl_readdata[10]~q ),
	.dma_ctl_readdata_11(\dma_1|dma_ctl_readdata[11]~q ),
	.dma_ctl_readdata_12(\dma_1|dma_ctl_readdata[12]~q ),
	.dma_ctl_readdata_13(\dma_1|dma_ctl_readdata[13]~q ),
	.dma_ctl_readdata_14(\dma_1|dma_ctl_readdata[14]~q ),
	.dma_ctl_readdata_15(\dma_1|dma_ctl_readdata[15]~q ),
	.dma_ctl_readdata_16(\dma_1|dma_ctl_readdata[16]~q ),
	.dma_ctl_readdata_17(\dma_1|dma_ctl_readdata[17]~q ),
	.dma_ctl_readdata_18(\dma_1|dma_ctl_readdata[18]~q ),
	.dma_ctl_readdata_19(\dma_1|dma_ctl_readdata[19]~q ),
	.dma_ctl_readdata_20(\dma_1|dma_ctl_readdata[20]~q ),
	.dma_ctl_readdata_21(\dma_1|dma_ctl_readdata[21]~q ),
	.dma_ctl_readdata_22(\dma_1|dma_ctl_readdata[22]~q ),
	.dma_ctl_readdata_23(\dma_1|dma_ctl_readdata[23]~q ),
	.dma_ctl_readdata_24(\dma_1|dma_ctl_readdata[24]~q ),
	.dma_ctl_readdata_25(\dma_1|dma_ctl_readdata[25]~q ),
	.dma_ctl_readdata_26(\dma_1|dma_ctl_readdata[26]~q ),
	.dma_ctl_readdata_27(\dma_1|dma_ctl_readdata[27]~q ),
	.dma_ctl_readdata_28(\dma_1|dma_ctl_readdata[28]~q ),
	.dma_ctl_readdata_29(\dma_1|dma_ctl_readdata[29]~q ),
	.dma_ctl_readdata_30(\dma_1|dma_ctl_readdata[30]~q ),
	.dma_ctl_readdata_31(\dma_1|dma_ctl_readdata[31]~q ),
	.av_readdatavalid4(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~4_combout ),
	.src0_valid(\mm_interconnect_1|rsp_demux|src0_valid~1_combout ),
	.src_data_8(\mm_interconnect_1|rsp_mux|src_data[8]~0_combout ),
	.src_data_81(\mm_interconnect_1|rsp_mux|src_data[8]~1_combout ),
	.src_data_16(\mm_interconnect_1|rsp_mux|src_data[16]~4_combout ),
	.src_data_24(\mm_interconnect_1|rsp_mux|src_data[24]~7_combout ),
	.src_data_0(\mm_interconnect_1|rsp_mux|src_data[0]~8_combout ),
	.src_data_01(\mm_interconnect_1|rsp_mux|src_data[0]~9_combout ),
	.in_data_reg_0(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_1(\mm_interconnect_0|dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.src_data_9(\mm_interconnect_1|rsp_mux|src_data[9]~10_combout ),
	.src_data_91(\mm_interconnect_1|rsp_mux|src_data[9]~11_combout ),
	.src_data_17(\mm_interconnect_1|rsp_mux|src_data[17]~14_combout ),
	.src_data_25(\mm_interconnect_1|rsp_mux|src_data[25]~17_combout ),
	.src_data_1(\mm_interconnect_1|rsp_mux|src_data[1]~18_combout ),
	.src_data_11(\mm_interconnect_1|rsp_mux|src_data[1]~19_combout ),
	.src_data_10(\mm_interconnect_1|rsp_mux|src_data[10]~20_combout ),
	.src_data_101(\mm_interconnect_1|rsp_mux|src_data[10]~21_combout ),
	.src_data_18(\mm_interconnect_1|rsp_mux|src_data[18]~24_combout ),
	.src_data_26(\mm_interconnect_1|rsp_mux|src_data[26]~27_combout ),
	.src_data_2(\mm_interconnect_1|rsp_mux|src_data[2]~28_combout ),
	.src_data_21(\mm_interconnect_1|rsp_mux|src_data[2]~29_combout ),
	.src_data_111(\mm_interconnect_1|rsp_mux|src_data[11]~30_combout ),
	.src_data_112(\mm_interconnect_1|rsp_mux|src_data[11]~31_combout ),
	.src_data_19(\mm_interconnect_1|rsp_mux|src_data[19]~34_combout ),
	.src_data_27(\mm_interconnect_1|rsp_mux|src_data[27]~37_combout ),
	.src_data_3(\mm_interconnect_1|rsp_mux|src_data[3]~38_combout ),
	.src_data_31(\mm_interconnect_1|rsp_mux|src_data[3]~39_combout ),
	.src_data_12(\mm_interconnect_1|rsp_mux|src_data[12]~40_combout ),
	.src_data_121(\mm_interconnect_1|rsp_mux|src_data[12]~41_combout ),
	.src_data_20(\mm_interconnect_1|rsp_mux|src_data[20]~44_combout ),
	.src_data_28(\mm_interconnect_1|rsp_mux|src_data[28]~47_combout ),
	.src_data_4(\mm_interconnect_1|rsp_mux|src_data[4]~48_combout ),
	.src_data_41(\mm_interconnect_1|rsp_mux|src_data[4]~49_combout ),
	.src_data_13(\mm_interconnect_1|rsp_mux|src_data[13]~50_combout ),
	.src_data_131(\mm_interconnect_1|rsp_mux|src_data[13]~51_combout ),
	.src_data_211(\mm_interconnect_1|rsp_mux|src_data[21]~54_combout ),
	.src_data_29(\mm_interconnect_1|rsp_mux|src_data[29]~57_combout ),
	.src_data_5(\mm_interconnect_1|rsp_mux|src_data[5]~58_combout ),
	.src_data_51(\mm_interconnect_1|rsp_mux|src_data[5]~59_combout ),
	.src_data_14(\mm_interconnect_1|rsp_mux|src_data[14]~60_combout ),
	.src_data_141(\mm_interconnect_1|rsp_mux|src_data[14]~61_combout ),
	.src_data_22(\mm_interconnect_1|rsp_mux|src_data[22]~64_combout ),
	.src_data_30(\mm_interconnect_1|rsp_mux|src_data[30]~67_combout ),
	.src_data_6(\mm_interconnect_1|rsp_mux|src_data[6]~68_combout ),
	.src_data_61(\mm_interconnect_1|rsp_mux|src_data[6]~69_combout ),
	.src_data_15(\mm_interconnect_1|rsp_mux|src_data[15]~70_combout ),
	.src_data_151(\mm_interconnect_1|rsp_mux|src_data[15]~71_combout ),
	.src_data_23(\mm_interconnect_1|rsp_mux|src_data[23]~74_combout ),
	.src_data_311(\mm_interconnect_1|rsp_mux|src_data[31]~77_combout ),
	.src_data_7(\mm_interconnect_1|rsp_mux|src_data[7]~78_combout ),
	.src_data_71(\mm_interconnect_1|rsp_mux|src_data[7]~79_combout ),
	.src_data_82(\mm_interconnect_1|rsp_mux|src_data[8]~80_combout ),
	.src_data_92(\mm_interconnect_1|rsp_mux|src_data[9]~81_combout ),
	.src_data_102(\mm_interconnect_1|rsp_mux|src_data[10]~82_combout ),
	.src_data_113(\mm_interconnect_1|rsp_mux|src_data[11]~83_combout ),
	.src_data_122(\mm_interconnect_1|rsp_mux|src_data[12]~84_combout ),
	.src_data_132(\mm_interconnect_1|rsp_mux|src_data[13]~85_combout ),
	.src_data_142(\mm_interconnect_1|rsp_mux|src_data[14]~86_combout ),
	.src_data_152(\mm_interconnect_1|rsp_mux|src_data[15]~87_combout ));

Computer_System_Computer_System_System_PLL system_pll(
	.outclk_wire_1(\system_pll|sys_pll|altera_pll_i|outclk_wire[1] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.locked_wire_0(\system_pll|sys_pll|altera_pll_i|locked_wire[0] ),
	.system_pll_ref_clk_clk(\system_pll_ref_clk_clk~input_o ),
	.system_pll_ref_reset_reset(\system_pll_ref_reset_reset~input_o ));

Computer_System_Computer_System_mm_interconnect_1 mm_interconnect_1(
	.f2h_ARREADY_0(\arm_a9_hps|fpga_interfaces|f2h_ARREADY[0] ),
	.f2h_AWREADY_0(\arm_a9_hps|fpga_interfaces|f2h_AWREADY[0] ),
	.f2h_BVALID_0(\arm_a9_hps|fpga_interfaces|f2h_BVALID[0] ),
	.f2h_RVALID_0(\arm_a9_hps|fpga_interfaces|f2h_RVALID[0] ),
	.f2h_WREADY_0(\arm_a9_hps|fpga_interfaces|f2h_WREADY[0] ),
	.f2h_RDATA_0(\arm_a9_hps|fpga_interfaces|f2h_RDATA[0] ),
	.f2h_RDATA_1(\arm_a9_hps|fpga_interfaces|f2h_RDATA[1] ),
	.f2h_RDATA_2(\arm_a9_hps|fpga_interfaces|f2h_RDATA[2] ),
	.f2h_RDATA_3(\arm_a9_hps|fpga_interfaces|f2h_RDATA[3] ),
	.f2h_RDATA_4(\arm_a9_hps|fpga_interfaces|f2h_RDATA[4] ),
	.f2h_RDATA_5(\arm_a9_hps|fpga_interfaces|f2h_RDATA[5] ),
	.f2h_RDATA_6(\arm_a9_hps|fpga_interfaces|f2h_RDATA[6] ),
	.f2h_RDATA_7(\arm_a9_hps|fpga_interfaces|f2h_RDATA[7] ),
	.f2h_RDATA_8(\arm_a9_hps|fpga_interfaces|f2h_RDATA[8] ),
	.f2h_RDATA_9(\arm_a9_hps|fpga_interfaces|f2h_RDATA[9] ),
	.f2h_RDATA_10(\arm_a9_hps|fpga_interfaces|f2h_RDATA[10] ),
	.f2h_RDATA_11(\arm_a9_hps|fpga_interfaces|f2h_RDATA[11] ),
	.f2h_RDATA_12(\arm_a9_hps|fpga_interfaces|f2h_RDATA[12] ),
	.f2h_RDATA_13(\arm_a9_hps|fpga_interfaces|f2h_RDATA[13] ),
	.f2h_RDATA_14(\arm_a9_hps|fpga_interfaces|f2h_RDATA[14] ),
	.f2h_RDATA_15(\arm_a9_hps|fpga_interfaces|f2h_RDATA[15] ),
	.f2h_RDATA_16(\arm_a9_hps|fpga_interfaces|f2h_RDATA[16] ),
	.f2h_RDATA_17(\arm_a9_hps|fpga_interfaces|f2h_RDATA[17] ),
	.f2h_RDATA_18(\arm_a9_hps|fpga_interfaces|f2h_RDATA[18] ),
	.f2h_RDATA_19(\arm_a9_hps|fpga_interfaces|f2h_RDATA[19] ),
	.f2h_RDATA_20(\arm_a9_hps|fpga_interfaces|f2h_RDATA[20] ),
	.f2h_RDATA_21(\arm_a9_hps|fpga_interfaces|f2h_RDATA[21] ),
	.f2h_RDATA_22(\arm_a9_hps|fpga_interfaces|f2h_RDATA[22] ),
	.f2h_RDATA_23(\arm_a9_hps|fpga_interfaces|f2h_RDATA[23] ),
	.f2h_RDATA_24(\arm_a9_hps|fpga_interfaces|f2h_RDATA[24] ),
	.f2h_RDATA_25(\arm_a9_hps|fpga_interfaces|f2h_RDATA[25] ),
	.f2h_RDATA_26(\arm_a9_hps|fpga_interfaces|f2h_RDATA[26] ),
	.f2h_RDATA_27(\arm_a9_hps|fpga_interfaces|f2h_RDATA[27] ),
	.f2h_RDATA_28(\arm_a9_hps|fpga_interfaces|f2h_RDATA[28] ),
	.f2h_RDATA_29(\arm_a9_hps|fpga_interfaces|f2h_RDATA[29] ),
	.f2h_RDATA_30(\arm_a9_hps|fpga_interfaces|f2h_RDATA[30] ),
	.f2h_RDATA_31(\arm_a9_hps|fpga_interfaces|f2h_RDATA[31] ),
	.f2h_RDATA_32(\arm_a9_hps|fpga_interfaces|f2h_RDATA[32] ),
	.f2h_RDATA_33(\arm_a9_hps|fpga_interfaces|f2h_RDATA[33] ),
	.f2h_RDATA_34(\arm_a9_hps|fpga_interfaces|f2h_RDATA[34] ),
	.f2h_RDATA_35(\arm_a9_hps|fpga_interfaces|f2h_RDATA[35] ),
	.f2h_RDATA_36(\arm_a9_hps|fpga_interfaces|f2h_RDATA[36] ),
	.f2h_RDATA_37(\arm_a9_hps|fpga_interfaces|f2h_RDATA[37] ),
	.f2h_RDATA_38(\arm_a9_hps|fpga_interfaces|f2h_RDATA[38] ),
	.f2h_RDATA_39(\arm_a9_hps|fpga_interfaces|f2h_RDATA[39] ),
	.f2h_RDATA_40(\arm_a9_hps|fpga_interfaces|f2h_RDATA[40] ),
	.f2h_RDATA_41(\arm_a9_hps|fpga_interfaces|f2h_RDATA[41] ),
	.f2h_RDATA_42(\arm_a9_hps|fpga_interfaces|f2h_RDATA[42] ),
	.f2h_RDATA_43(\arm_a9_hps|fpga_interfaces|f2h_RDATA[43] ),
	.f2h_RDATA_44(\arm_a9_hps|fpga_interfaces|f2h_RDATA[44] ),
	.f2h_RDATA_45(\arm_a9_hps|fpga_interfaces|f2h_RDATA[45] ),
	.f2h_RDATA_46(\arm_a9_hps|fpga_interfaces|f2h_RDATA[46] ),
	.f2h_RDATA_47(\arm_a9_hps|fpga_interfaces|f2h_RDATA[47] ),
	.f2h_RDATA_48(\arm_a9_hps|fpga_interfaces|f2h_RDATA[48] ),
	.f2h_RDATA_49(\arm_a9_hps|fpga_interfaces|f2h_RDATA[49] ),
	.f2h_RDATA_50(\arm_a9_hps|fpga_interfaces|f2h_RDATA[50] ),
	.f2h_RDATA_51(\arm_a9_hps|fpga_interfaces|f2h_RDATA[51] ),
	.f2h_RDATA_52(\arm_a9_hps|fpga_interfaces|f2h_RDATA[52] ),
	.f2h_RDATA_53(\arm_a9_hps|fpga_interfaces|f2h_RDATA[53] ),
	.f2h_RDATA_54(\arm_a9_hps|fpga_interfaces|f2h_RDATA[54] ),
	.f2h_RDATA_55(\arm_a9_hps|fpga_interfaces|f2h_RDATA[55] ),
	.f2h_RDATA_56(\arm_a9_hps|fpga_interfaces|f2h_RDATA[56] ),
	.f2h_RDATA_57(\arm_a9_hps|fpga_interfaces|f2h_RDATA[57] ),
	.f2h_RDATA_58(\arm_a9_hps|fpga_interfaces|f2h_RDATA[58] ),
	.f2h_RDATA_59(\arm_a9_hps|fpga_interfaces|f2h_RDATA[59] ),
	.f2h_RDATA_60(\arm_a9_hps|fpga_interfaces|f2h_RDATA[60] ),
	.f2h_RDATA_61(\arm_a9_hps|fpga_interfaces|f2h_RDATA[61] ),
	.f2h_RDATA_62(\arm_a9_hps|fpga_interfaces|f2h_RDATA[62] ),
	.f2h_RDATA_63(\arm_a9_hps|fpga_interfaces|f2h_RDATA[63] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.readaddress_2(\dma_1|readaddress[2]~q ),
	.readaddress_3(\dma_1|readaddress[3]~q ),
	.readaddress_4(\dma_1|readaddress[4]~q ),
	.readaddress_5(\dma_1|readaddress[5]~q ),
	.readaddress_6(\dma_1|readaddress[6]~q ),
	.readaddress_7(\dma_1|readaddress[7]~q ),
	.readaddress_8(\dma_1|readaddress[8]~q ),
	.readaddress_9(\dma_1|readaddress[9]~q ),
	.readaddress_10(\dma_1|readaddress[10]~q ),
	.readaddress_11(\dma_1|readaddress[11]~q ),
	.readaddress_12(\dma_1|readaddress[12]~q ),
	.readaddress_13(\dma_1|readaddress[13]~q ),
	.readaddress_14(\dma_1|readaddress[14]~q ),
	.readaddress_15(\dma_1|readaddress[15]~q ),
	.readaddress_16(\dma_1|readaddress[16]~q ),
	.readaddress_17(\dma_1|readaddress[17]~q ),
	.readaddress_18(\dma_1|readaddress[18]~q ),
	.readaddress_19(\dma_1|readaddress[19]~q ),
	.readaddress_20(\dma_1|readaddress[20]~q ),
	.readaddress_21(\dma_1|readaddress[21]~q ),
	.readaddress_22(\dma_1|readaddress[22]~q ),
	.readaddress_23(\dma_1|readaddress[23]~q ),
	.readaddress_24(\dma_1|readaddress[24]~q ),
	.readaddress_25(\dma_1|readaddress[25]~q ),
	.readaddress_26(\dma_1|readaddress[26]~q ),
	.readaddress_27(\dma_1|readaddress[27]~q ),
	.readaddress_28(\dma_1|readaddress[28]~q ),
	.readaddress_29(\dma_1|readaddress[29]~q ),
	.readaddress_30(\dma_1|readaddress[30]~q ),
	.readaddress_31(\dma_1|readaddress[31]~q ),
	.writeaddress_2(\dma_2|writeaddress[2]~q ),
	.writeaddress_3(\dma_2|writeaddress[3]~q ),
	.writeaddress_4(\dma_2|writeaddress[4]~q ),
	.writeaddress_5(\dma_2|writeaddress[5]~q ),
	.writeaddress_6(\dma_2|writeaddress[6]~q ),
	.writeaddress_7(\dma_2|writeaddress[7]~q ),
	.writeaddress_8(\dma_2|writeaddress[8]~q ),
	.writeaddress_9(\dma_2|writeaddress[9]~q ),
	.writeaddress_10(\dma_2|writeaddress[10]~q ),
	.writeaddress_11(\dma_2|writeaddress[11]~q ),
	.writeaddress_12(\dma_2|writeaddress[12]~q ),
	.writeaddress_13(\dma_2|writeaddress[13]~q ),
	.writeaddress_14(\dma_2|writeaddress[14]~q ),
	.writeaddress_15(\dma_2|writeaddress[15]~q ),
	.writeaddress_16(\dma_2|writeaddress[16]~q ),
	.writeaddress_17(\dma_2|writeaddress[17]~q ),
	.writeaddress_18(\dma_2|writeaddress[18]~q ),
	.writeaddress_19(\dma_2|writeaddress[19]~q ),
	.writeaddress_20(\dma_2|writeaddress[20]~q ),
	.writeaddress_21(\dma_2|writeaddress[21]~q ),
	.writeaddress_22(\dma_2|writeaddress[22]~q ),
	.writeaddress_23(\dma_2|writeaddress[23]~q ),
	.writeaddress_24(\dma_2|writeaddress[24]~q ),
	.writeaddress_25(\dma_2|writeaddress[25]~q ),
	.writeaddress_26(\dma_2|writeaddress[26]~q ),
	.writeaddress_27(\dma_2|writeaddress[27]~q ),
	.writeaddress_28(\dma_2|writeaddress[28]~q ),
	.writeaddress_29(\dma_2|writeaddress[29]~q ),
	.writeaddress_30(\dma_2|writeaddress[30]~q ),
	.writeaddress_31(\dma_2|writeaddress[31]~q ),
	.q_b_0(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[0] ),
	.q_b_1(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[1] ),
	.q_b_2(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[2] ),
	.q_b_3(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[3] ),
	.q_b_4(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[4] ),
	.q_b_5(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[5] ),
	.q_b_6(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[6] ),
	.q_b_7(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[7] ),
	.q_b_8(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[8] ),
	.q_b_9(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[9] ),
	.q_b_10(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[10] ),
	.q_b_11(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[11] ),
	.q_b_12(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[12] ),
	.q_b_13(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[13] ),
	.q_b_14(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[14] ),
	.q_b_15(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[15] ),
	.q_b_16(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[16] ),
	.q_b_17(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[17] ),
	.q_b_18(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[18] ),
	.q_b_19(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[19] ),
	.q_b_20(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[20] ),
	.q_b_21(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[21] ),
	.q_b_22(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[22] ),
	.q_b_23(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[23] ),
	.q_b_24(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[24] ),
	.q_b_25(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[25] ),
	.q_b_26(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[26] ),
	.q_b_27(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[27] ),
	.q_b_28(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[28] ),
	.q_b_29(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[29] ),
	.q_b_30(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[30] ),
	.q_b_31(\dma_2|the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[31] ),
	.writeaddress_1(\dma_2|writeaddress[1]~q ),
	.writeaddress_0(\dma_2|writeaddress[0]~q ),
	.mem_used_7(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem_used[7]~q ),
	.saved_grant_0(\mm_interconnect_1|cmd_mux_001|saved_grant[0]~q ),
	.read_select(\dma_1|the_Computer_System_dma_1_mem_read|read_select~q ),
	.hold_waitrequest(\mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ),
	.write(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|write~0_combout ),
	.arvalid(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|arvalid~combout ),
	.address_taken(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|address_taken~q ),
	.mem_used_71(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[7]~q ),
	.fifo_empty(\dma_2|the_Computer_System_dma_2_fifo_module|fifo_empty~q ),
	.saved_grant_1(\mm_interconnect_1|cmd_mux|saved_grant[1]~q ),
	.src_valid(\mm_interconnect_1|cmd_mux|src_valid~0_combout ),
	.awvalid(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|awvalid~combout ),
	.ARM_A9_HPS_f2h_axi_slave_bready(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|bready~0_combout ),
	.data_taken(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|data_taken~q ),
	.wvalid(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|wvalid~combout ),
	.src_payload(\mm_interconnect_1|cmd_mux_001|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_1|cmd_mux_001|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_1|cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_1|cmd_mux_001|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_1|cmd_mux_001|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_1|cmd_mux_001|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_1|cmd_mux_001|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_1|cmd_mux_001|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_1|cmd_mux_001|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_1|cmd_mux_001|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_1|cmd_mux_001|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_1|cmd_mux_001|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_1|cmd_mux_001|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_1|cmd_mux_001|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_1|cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_1|cmd_mux_001|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_1|cmd_mux_001|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_1|cmd_mux_001|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_1|cmd_mux_001|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_1|cmd_mux_001|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_1|cmd_mux_001|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_1|cmd_mux_001|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_1|cmd_mux_001|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_1|cmd_mux_001|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_1|cmd_mux_001|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_1|cmd_mux_001|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_1|cmd_mux_001|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_1|cmd_mux_001|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_1|cmd_mux_001|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_1|cmd_mux_001|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_1|cmd_mux|src_payload~0_combout ),
	.src_payload31(\mm_interconnect_1|cmd_mux|src_payload~1_combout ),
	.src_payload32(\mm_interconnect_1|cmd_mux|src_payload~2_combout ),
	.src_payload33(\mm_interconnect_1|cmd_mux|src_payload~3_combout ),
	.src_payload34(\mm_interconnect_1|cmd_mux|src_payload~4_combout ),
	.src_payload35(\mm_interconnect_1|cmd_mux|src_payload~5_combout ),
	.src_payload36(\mm_interconnect_1|cmd_mux|src_payload~6_combout ),
	.src_payload37(\mm_interconnect_1|cmd_mux|src_payload~7_combout ),
	.src_payload38(\mm_interconnect_1|cmd_mux|src_payload~8_combout ),
	.src_payload39(\mm_interconnect_1|cmd_mux|src_payload~9_combout ),
	.src_payload40(\mm_interconnect_1|cmd_mux|src_payload~10_combout ),
	.src_payload41(\mm_interconnect_1|cmd_mux|src_payload~11_combout ),
	.src_payload42(\mm_interconnect_1|cmd_mux|src_payload~12_combout ),
	.src_payload43(\mm_interconnect_1|cmd_mux|src_payload~13_combout ),
	.src_payload44(\mm_interconnect_1|cmd_mux|src_payload~14_combout ),
	.src_payload45(\mm_interconnect_1|cmd_mux|src_payload~15_combout ),
	.src_payload46(\mm_interconnect_1|cmd_mux|src_payload~16_combout ),
	.src_payload47(\mm_interconnect_1|cmd_mux|src_payload~17_combout ),
	.src_payload48(\mm_interconnect_1|cmd_mux|src_payload~18_combout ),
	.src_payload49(\mm_interconnect_1|cmd_mux|src_payload~19_combout ),
	.src_payload50(\mm_interconnect_1|cmd_mux|src_payload~20_combout ),
	.src_payload51(\mm_interconnect_1|cmd_mux|src_payload~21_combout ),
	.src_payload52(\mm_interconnect_1|cmd_mux|src_payload~22_combout ),
	.src_payload53(\mm_interconnect_1|cmd_mux|src_payload~23_combout ),
	.src_payload54(\mm_interconnect_1|cmd_mux|src_payload~24_combout ),
	.src_payload55(\mm_interconnect_1|cmd_mux|src_payload~25_combout ),
	.src_payload56(\mm_interconnect_1|cmd_mux|src_payload~26_combout ),
	.src_payload57(\mm_interconnect_1|cmd_mux|src_payload~27_combout ),
	.src_payload58(\mm_interconnect_1|cmd_mux|src_payload~28_combout ),
	.src_payload59(\mm_interconnect_1|cmd_mux|src_payload~29_combout ),
	.last_write_collision(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_collision~q ),
	.last_write_data_0(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[0]~q ),
	.control_2(\dma_2|control[2]~q ),
	.control_0(\dma_2|control[0]~q ),
	.ShiftLeft1(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~0_combout ),
	.last_write_data_1(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[1]~q ),
	.ShiftLeft11(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~1_combout ),
	.last_write_data_2(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[2]~q ),
	.ShiftLeft12(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~2_combout ),
	.last_write_data_3(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[3]~q ),
	.ShiftLeft13(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~3_combout ),
	.last_write_data_4(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[4]~q ),
	.ShiftLeft14(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~4_combout ),
	.last_write_data_5(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[5]~q ),
	.ShiftLeft15(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~5_combout ),
	.last_write_data_6(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[6]~q ),
	.ShiftLeft16(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~6_combout ),
	.last_write_data_7(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[7]~q ),
	.ShiftLeft17(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~7_combout ),
	.write_writedata(\dma_2|write_writedata~0_combout ),
	.last_write_data_8(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[8]~q ),
	.ShiftLeft18(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~9_combout ),
	.write_writedata1(\dma_2|write_writedata~1_combout ),
	.last_write_data_9(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[9]~q ),
	.ShiftLeft19(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~11_combout ),
	.write_writedata2(\dma_2|write_writedata~2_combout ),
	.last_write_data_10(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[10]~q ),
	.ShiftLeft110(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~13_combout ),
	.write_writedata3(\dma_2|write_writedata~3_combout ),
	.last_write_data_11(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[11]~q ),
	.ShiftLeft111(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~15_combout ),
	.write_writedata4(\dma_2|write_writedata~4_combout ),
	.last_write_data_12(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[12]~q ),
	.ShiftLeft112(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~17_combout ),
	.write_writedata5(\dma_2|write_writedata~5_combout ),
	.last_write_data_13(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[13]~q ),
	.ShiftLeft113(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~19_combout ),
	.write_writedata6(\dma_2|write_writedata~6_combout ),
	.last_write_data_14(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[14]~q ),
	.ShiftLeft114(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~21_combout ),
	.write_writedata7(\dma_2|write_writedata~7_combout ),
	.last_write_data_15(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[15]~q ),
	.ShiftLeft115(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~23_combout ),
	.last_write_data_16(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[16]~q ),
	.ShiftLeft116(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~25_combout ),
	.last_write_data_17(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[17]~q ),
	.ShiftLeft117(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~27_combout ),
	.last_write_data_18(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[18]~q ),
	.ShiftLeft118(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~29_combout ),
	.last_write_data_19(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[19]~q ),
	.ShiftLeft119(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~31_combout ),
	.last_write_data_20(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[20]~q ),
	.ShiftLeft120(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~33_combout ),
	.last_write_data_21(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[21]~q ),
	.ShiftLeft121(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~35_combout ),
	.last_write_data_22(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[22]~q ),
	.ShiftLeft122(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~37_combout ),
	.last_write_data_23(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[23]~q ),
	.ShiftLeft123(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~39_combout ),
	.last_write_data_24(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[24]~q ),
	.ShiftLeft124(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~41_combout ),
	.last_write_data_25(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[25]~q ),
	.ShiftLeft125(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~43_combout ),
	.last_write_data_26(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[26]~q ),
	.ShiftLeft126(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~45_combout ),
	.last_write_data_27(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[27]~q ),
	.ShiftLeft127(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~47_combout ),
	.last_write_data_28(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[28]~q ),
	.ShiftLeft128(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~49_combout ),
	.last_write_data_29(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[29]~q ),
	.ShiftLeft129(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~51_combout ),
	.last_write_data_30(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[30]~q ),
	.ShiftLeft130(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~53_combout ),
	.last_write_data_31(\dma_2|the_Computer_System_dma_2_fifo_module|last_write_data[31]~q ),
	.ShiftLeft131(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~55_combout ),
	.ShiftLeft132(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~56_combout ),
	.ShiftLeft133(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~57_combout ),
	.ShiftLeft134(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~58_combout ),
	.ShiftLeft135(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~59_combout ),
	.ShiftLeft136(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~60_combout ),
	.ShiftLeft137(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~61_combout ),
	.ShiftLeft138(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~62_combout ),
	.ShiftLeft139(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~63_combout ),
	.ShiftLeft140(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~64_combout ),
	.ShiftLeft141(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~65_combout ),
	.ShiftLeft142(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~66_combout ),
	.ShiftLeft143(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~67_combout ),
	.ShiftLeft144(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~68_combout ),
	.ShiftLeft145(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~69_combout ),
	.ShiftLeft146(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~70_combout ),
	.ShiftLeft147(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~71_combout ),
	.ShiftLeft148(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~72_combout ),
	.ShiftLeft149(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~73_combout ),
	.ShiftLeft150(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~74_combout ),
	.ShiftLeft151(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~75_combout ),
	.ShiftLeft152(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~76_combout ),
	.ShiftLeft153(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~77_combout ),
	.ShiftLeft154(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~78_combout ),
	.ShiftLeft155(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~79_combout ),
	.ShiftLeft156(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~80_combout ),
	.ShiftLeft157(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~81_combout ),
	.ShiftLeft158(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~82_combout ),
	.ShiftLeft159(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~83_combout ),
	.ShiftLeft160(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~84_combout ),
	.ShiftLeft161(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~85_combout ),
	.ShiftLeft162(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~86_combout ),
	.ShiftLeft163(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft1~87_combout ),
	.ShiftLeft0(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~0_combout ),
	.ShiftLeft01(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~1_combout ),
	.ShiftLeft02(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~2_combout ),
	.ShiftLeft03(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~3_combout ),
	.ShiftLeft04(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~4_combout ),
	.ShiftLeft05(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~5_combout ),
	.ShiftLeft06(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~6_combout ),
	.ShiftLeft07(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter|ShiftLeft0~7_combout ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.WideOr1(\mm_interconnect_1|cmd_mux_001|WideOr1~0_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.inc_read(\dma_1|the_Computer_System_dma_1_mem_read|inc_read~combout ),
	.av_readdatavalid(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~0_combout ),
	.av_readdatavalid1(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~1_combout ),
	.av_readdatavalid2(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~2_combout ),
	.av_readdatavalid3(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~3_combout ),
	.fifo_read(\dma_2|the_Computer_System_dma_2_mem_write|fifo_read~0_combout ),
	.write_cp_ready(\mm_interconnect_1|arm_a9_hps_f2h_axi_slave_agent|write_cp_ready~0_combout ),
	.av_readdatavalid4(\mm_interconnect_1|dma_1_read_master_agent|av_readdatavalid~4_combout ),
	.src0_valid(\mm_interconnect_1|rsp_demux|src0_valid~1_combout ),
	.src_data_8(\mm_interconnect_1|rsp_mux|src_data[8]~0_combout ),
	.src_data_81(\mm_interconnect_1|rsp_mux|src_data[8]~1_combout ),
	.src_data_16(\mm_interconnect_1|rsp_mux|src_data[16]~4_combout ),
	.src_data_24(\mm_interconnect_1|rsp_mux|src_data[24]~7_combout ),
	.src_data_0(\mm_interconnect_1|rsp_mux|src_data[0]~8_combout ),
	.src_data_01(\mm_interconnect_1|rsp_mux|src_data[0]~9_combout ),
	.src_data_9(\mm_interconnect_1|rsp_mux|src_data[9]~10_combout ),
	.src_data_91(\mm_interconnect_1|rsp_mux|src_data[9]~11_combout ),
	.src_data_17(\mm_interconnect_1|rsp_mux|src_data[17]~14_combout ),
	.src_data_25(\mm_interconnect_1|rsp_mux|src_data[25]~17_combout ),
	.src_data_1(\mm_interconnect_1|rsp_mux|src_data[1]~18_combout ),
	.src_data_11(\mm_interconnect_1|rsp_mux|src_data[1]~19_combout ),
	.src_data_10(\mm_interconnect_1|rsp_mux|src_data[10]~20_combout ),
	.src_data_101(\mm_interconnect_1|rsp_mux|src_data[10]~21_combout ),
	.src_data_18(\mm_interconnect_1|rsp_mux|src_data[18]~24_combout ),
	.src_data_26(\mm_interconnect_1|rsp_mux|src_data[26]~27_combout ),
	.src_data_2(\mm_interconnect_1|rsp_mux|src_data[2]~28_combout ),
	.src_data_21(\mm_interconnect_1|rsp_mux|src_data[2]~29_combout ),
	.src_data_111(\mm_interconnect_1|rsp_mux|src_data[11]~30_combout ),
	.src_data_112(\mm_interconnect_1|rsp_mux|src_data[11]~31_combout ),
	.src_data_19(\mm_interconnect_1|rsp_mux|src_data[19]~34_combout ),
	.src_data_27(\mm_interconnect_1|rsp_mux|src_data[27]~37_combout ),
	.src_data_3(\mm_interconnect_1|rsp_mux|src_data[3]~38_combout ),
	.src_data_31(\mm_interconnect_1|rsp_mux|src_data[3]~39_combout ),
	.src_data_12(\mm_interconnect_1|rsp_mux|src_data[12]~40_combout ),
	.src_data_121(\mm_interconnect_1|rsp_mux|src_data[12]~41_combout ),
	.src_data_20(\mm_interconnect_1|rsp_mux|src_data[20]~44_combout ),
	.src_data_28(\mm_interconnect_1|rsp_mux|src_data[28]~47_combout ),
	.src_data_4(\mm_interconnect_1|rsp_mux|src_data[4]~48_combout ),
	.src_data_41(\mm_interconnect_1|rsp_mux|src_data[4]~49_combout ),
	.src_data_13(\mm_interconnect_1|rsp_mux|src_data[13]~50_combout ),
	.src_data_131(\mm_interconnect_1|rsp_mux|src_data[13]~51_combout ),
	.src_data_211(\mm_interconnect_1|rsp_mux|src_data[21]~54_combout ),
	.src_data_29(\mm_interconnect_1|rsp_mux|src_data[29]~57_combout ),
	.src_data_5(\mm_interconnect_1|rsp_mux|src_data[5]~58_combout ),
	.src_data_51(\mm_interconnect_1|rsp_mux|src_data[5]~59_combout ),
	.src_data_14(\mm_interconnect_1|rsp_mux|src_data[14]~60_combout ),
	.src_data_141(\mm_interconnect_1|rsp_mux|src_data[14]~61_combout ),
	.src_data_22(\mm_interconnect_1|rsp_mux|src_data[22]~64_combout ),
	.src_data_30(\mm_interconnect_1|rsp_mux|src_data[30]~67_combout ),
	.src_data_6(\mm_interconnect_1|rsp_mux|src_data[6]~68_combout ),
	.src_data_61(\mm_interconnect_1|rsp_mux|src_data[6]~69_combout ),
	.src_data_15(\mm_interconnect_1|rsp_mux|src_data[15]~70_combout ),
	.src_data_151(\mm_interconnect_1|rsp_mux|src_data[15]~71_combout ),
	.src_data_23(\mm_interconnect_1|rsp_mux|src_data[23]~74_combout ),
	.src_data_311(\mm_interconnect_1|rsp_mux|src_data[31]~77_combout ),
	.src_data_7(\mm_interconnect_1|rsp_mux|src_data[7]~78_combout ),
	.src_data_71(\mm_interconnect_1|rsp_mux|src_data[7]~79_combout ),
	.src_data_82(\mm_interconnect_1|rsp_mux|src_data[8]~80_combout ),
	.src_data_92(\mm_interconnect_1|rsp_mux|src_data[9]~81_combout ),
	.src_data_102(\mm_interconnect_1|rsp_mux|src_data[10]~82_combout ),
	.src_data_113(\mm_interconnect_1|rsp_mux|src_data[11]~83_combout ),
	.src_data_122(\mm_interconnect_1|rsp_mux|src_data[12]~84_combout ),
	.src_data_132(\mm_interconnect_1|rsp_mux|src_data[13]~85_combout ),
	.src_data_142(\mm_interconnect_1|rsp_mux|src_data[14]~86_combout ),
	.src_data_152(\mm_interconnect_1|rsp_mux|src_data[15]~87_combout ));

Computer_System_altera_reset_controller_1 rst_controller_001(
	.h2f_rst_n_0(\arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

Computer_System_altera_reset_controller rst_controller(
	.h2f_rst_n_0(\arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.locked_wire_0(\system_pll|sys_pll|altera_pll_i|locked_wire[0] ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.r_sync_rst1(\rst_controller|r_sync_rst~q ));

Computer_System_Computer_System_mm_interconnect_2 mm_interconnect_2(
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.readaddress_15(\dma_2|readaddress[15]~q ),
	.writeaddress_15(\dma_1|writeaddress[15]~q ),
	.q_b_0(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[0] ),
	.readaddress_2(\dma_2|readaddress[2]~q ),
	.writeaddress_2(\dma_1|writeaddress[2]~q ),
	.readaddress_3(\dma_2|readaddress[3]~q ),
	.writeaddress_3(\dma_1|writeaddress[3]~q ),
	.readaddress_4(\dma_2|readaddress[4]~q ),
	.writeaddress_4(\dma_1|writeaddress[4]~q ),
	.readaddress_5(\dma_2|readaddress[5]~q ),
	.writeaddress_5(\dma_1|writeaddress[5]~q ),
	.readaddress_6(\dma_2|readaddress[6]~q ),
	.writeaddress_6(\dma_1|writeaddress[6]~q ),
	.readaddress_7(\dma_2|readaddress[7]~q ),
	.writeaddress_7(\dma_1|writeaddress[7]~q ),
	.readaddress_8(\dma_2|readaddress[8]~q ),
	.writeaddress_8(\dma_1|writeaddress[8]~q ),
	.readaddress_9(\dma_2|readaddress[9]~q ),
	.writeaddress_9(\dma_1|writeaddress[9]~q ),
	.readaddress_10(\dma_2|readaddress[10]~q ),
	.writeaddress_10(\dma_1|writeaddress[10]~q ),
	.readaddress_11(\dma_2|readaddress[11]~q ),
	.writeaddress_11(\dma_1|writeaddress[11]~q ),
	.readaddress_12(\dma_2|readaddress[12]~q ),
	.writeaddress_12(\dma_1|writeaddress[12]~q ),
	.readaddress_13(\dma_2|readaddress[13]~q ),
	.writeaddress_13(\dma_1|writeaddress[13]~q ),
	.readaddress_14(\dma_2|readaddress[14]~q ),
	.writeaddress_14(\dma_1|writeaddress[14]~q ),
	.writeaddress_1(\dma_1|writeaddress[1]~q ),
	.writeaddress_0(\dma_1|writeaddress[0]~q ),
	.q_b_1(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[1] ),
	.q_b_2(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[2] ),
	.q_b_3(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[3] ),
	.q_b_4(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[4] ),
	.q_b_5(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[5] ),
	.q_b_6(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[6] ),
	.q_b_7(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[7] ),
	.q_b_8(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[8] ),
	.q_b_9(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[9] ),
	.q_b_10(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[10] ),
	.q_b_11(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[11] ),
	.q_b_12(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[12] ),
	.q_b_13(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[13] ),
	.q_b_14(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[14] ),
	.q_b_15(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[15] ),
	.q_b_16(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[16] ),
	.q_b_17(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[17] ),
	.q_b_18(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[18] ),
	.q_b_19(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[19] ),
	.q_b_20(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[20] ),
	.q_b_21(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[21] ),
	.q_b_22(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[22] ),
	.q_b_23(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[23] ),
	.q_b_24(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[24] ),
	.q_b_25(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[25] ),
	.q_b_26(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[26] ),
	.q_b_27(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[27] ),
	.q_b_28(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[28] ),
	.q_b_29(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[29] ),
	.q_b_30(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[30] ),
	.q_b_31(\dma_1|the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp_component|sram|ram_block|auto_generated|q_b[31] ),
	.hold_waitrequest(\mm_interconnect_2|dma_1_write_master_agent|hold_waitrequest~q ),
	.saved_grant_0(\mm_interconnect_2|cmd_mux|saved_grant[0]~q ),
	.saved_grant_1(\mm_interconnect_2|cmd_mux|saved_grant[1]~q ),
	.mem_used_1(\mm_interconnect_2|onchip_sram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.fifo_empty(\dma_1|the_Computer_System_dma_1_fifo_module|fifo_empty~q ),
	.last_write_collision(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_collision~q ),
	.last_write_data_0(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[0]~q ),
	.control_2(\dma_1|control[2]~q ),
	.control_0(\dma_1|control[0]~q ),
	.src_payload(\mm_interconnect_2|cmd_mux|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_2|cmd_mux|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_2|cmd_mux|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_2|cmd_mux|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_2|cmd_mux|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_2|cmd_mux|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_2|cmd_mux|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_2|cmd_mux|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_2|cmd_mux|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_2|cmd_mux|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_2|cmd_mux|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_2|cmd_mux|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_2|cmd_mux|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_2|cmd_mux|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_2|cmd_mux|src_data[32]~0_combout ),
	.last_write_data_1(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[1]~q ),
	.src_payload1(\mm_interconnect_2|cmd_mux|src_payload~2_combout ),
	.last_write_data_2(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[2]~q ),
	.src_payload2(\mm_interconnect_2|cmd_mux|src_payload~3_combout ),
	.last_write_data_3(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[3]~q ),
	.src_payload3(\mm_interconnect_2|cmd_mux|src_payload~4_combout ),
	.last_write_data_4(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[4]~q ),
	.src_payload4(\mm_interconnect_2|cmd_mux|src_payload~5_combout ),
	.last_write_data_5(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[5]~q ),
	.src_payload5(\mm_interconnect_2|cmd_mux|src_payload~6_combout ),
	.last_write_data_6(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[6]~q ),
	.src_payload6(\mm_interconnect_2|cmd_mux|src_payload~7_combout ),
	.last_write_data_7(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[7]~q ),
	.src_payload7(\mm_interconnect_2|cmd_mux|src_payload~8_combout ),
	.write_writedata(\dma_1|write_writedata~0_combout ),
	.last_write_data_8(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[8]~q ),
	.src_payload8(\mm_interconnect_2|cmd_mux|src_payload~9_combout ),
	.src_data_33(\mm_interconnect_2|cmd_mux|src_data[33]~1_combout ),
	.write_writedata1(\dma_1|write_writedata~1_combout ),
	.last_write_data_9(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[9]~q ),
	.src_payload9(\mm_interconnect_2|cmd_mux|src_payload~10_combout ),
	.write_writedata2(\dma_1|write_writedata~2_combout ),
	.last_write_data_10(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[10]~q ),
	.src_payload10(\mm_interconnect_2|cmd_mux|src_payload~11_combout ),
	.write_writedata3(\dma_1|write_writedata~3_combout ),
	.last_write_data_11(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[11]~q ),
	.src_payload11(\mm_interconnect_2|cmd_mux|src_payload~12_combout ),
	.write_writedata4(\dma_1|write_writedata~4_combout ),
	.last_write_data_12(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[12]~q ),
	.src_payload12(\mm_interconnect_2|cmd_mux|src_payload~13_combout ),
	.write_writedata5(\dma_1|write_writedata~5_combout ),
	.last_write_data_13(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[13]~q ),
	.src_payload13(\mm_interconnect_2|cmd_mux|src_payload~14_combout ),
	.write_writedata6(\dma_1|write_writedata~6_combout ),
	.last_write_data_14(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[14]~q ),
	.src_payload14(\mm_interconnect_2|cmd_mux|src_payload~15_combout ),
	.write_writedata7(\dma_1|write_writedata~7_combout ),
	.last_write_data_15(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[15]~q ),
	.src_payload15(\mm_interconnect_2|cmd_mux|src_payload~16_combout ),
	.last_write_data_16(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[16]~q ),
	.src_payload16(\mm_interconnect_2|cmd_mux|src_payload~17_combout ),
	.src_data_34(\mm_interconnect_2|cmd_mux|src_data[34]~2_combout ),
	.last_write_data_17(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[17]~q ),
	.src_payload17(\mm_interconnect_2|cmd_mux|src_payload~18_combout ),
	.last_write_data_18(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[18]~q ),
	.src_payload18(\mm_interconnect_2|cmd_mux|src_payload~19_combout ),
	.last_write_data_19(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[19]~q ),
	.src_payload19(\mm_interconnect_2|cmd_mux|src_payload~20_combout ),
	.last_write_data_20(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[20]~q ),
	.src_payload20(\mm_interconnect_2|cmd_mux|src_payload~21_combout ),
	.last_write_data_21(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[21]~q ),
	.src_payload21(\mm_interconnect_2|cmd_mux|src_payload~22_combout ),
	.last_write_data_22(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[22]~q ),
	.src_payload22(\mm_interconnect_2|cmd_mux|src_payload~23_combout ),
	.last_write_data_23(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[23]~q ),
	.src_payload23(\mm_interconnect_2|cmd_mux|src_payload~24_combout ),
	.last_write_data_24(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[24]~q ),
	.src_payload24(\mm_interconnect_2|cmd_mux|src_payload~25_combout ),
	.src_data_35(\mm_interconnect_2|cmd_mux|src_data[35]~3_combout ),
	.last_write_data_25(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[25]~q ),
	.src_payload25(\mm_interconnect_2|cmd_mux|src_payload~26_combout ),
	.last_write_data_26(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[26]~q ),
	.src_payload26(\mm_interconnect_2|cmd_mux|src_payload~27_combout ),
	.last_write_data_27(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[27]~q ),
	.src_payload27(\mm_interconnect_2|cmd_mux|src_payload~28_combout ),
	.last_write_data_28(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[28]~q ),
	.src_payload28(\mm_interconnect_2|cmd_mux|src_payload~29_combout ),
	.last_write_data_29(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[29]~q ),
	.src_payload29(\mm_interconnect_2|cmd_mux|src_payload~30_combout ),
	.last_write_data_30(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[30]~q ),
	.src_payload30(\mm_interconnect_2|cmd_mux|src_payload~31_combout ),
	.last_write_data_31(\dma_1|the_Computer_System_dma_1_fifo_module|last_write_data[31]~q ),
	.src_payload31(\mm_interconnect_2|cmd_mux|src_payload~32_combout ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.src0_valid(\mm_interconnect_2|rsp_demux|src0_valid~combout ),
	.read_select(\dma_2|the_Computer_System_dma_2_mem_read|read_select~q ),
	.read_latency_shift_reg(\mm_interconnect_2|onchip_sram_s1_translator|read_latency_shift_reg~0_combout ),
	.src_data_51(\mm_interconnect_2|cmd_mux|src_data[51]~combout ));

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[3]),
	.ibar(memory_mem_dqs_n[3]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[24]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[25]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[26]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[27]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[28]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[29]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[30]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[31]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[2]),
	.ibar(memory_mem_dqs_n[2]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[16]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[17]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[18]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[19]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[20]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[21]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[22]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[23]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[1]),
	.ibar(memory_mem_dqs_n[1]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[8]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[9]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[10]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[11]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[12]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[13]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[14]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[15]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[0]),
	.ibar(memory_mem_dqs_n[0]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[0]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[1]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[2]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[3]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[4]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[5]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[6]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[7]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

assign \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o  = hps_io_hps_io_emac1_inst_MDIO;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o  = hps_io_hps_io_qspi_inst_IO0;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o  = hps_io_hps_io_qspi_inst_IO1;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o  = hps_io_hps_io_qspi_inst_IO2;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o  = hps_io_hps_io_qspi_inst_IO3;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o  = hps_io_hps_io_sdio_inst_CMD;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o  = hps_io_hps_io_sdio_inst_D0;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o  = hps_io_hps_io_sdio_inst_D1;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o  = hps_io_hps_io_sdio_inst_D2;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o  = hps_io_hps_io_sdio_inst_D3;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~input_o  = hps_io_hps_io_usb1_inst_D0;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~input_o  = hps_io_hps_io_usb1_inst_D1;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~input_o  = hps_io_hps_io_usb1_inst_D2;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~input_o  = hps_io_hps_io_usb1_inst_D3;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~input_o  = hps_io_hps_io_usb1_inst_D4;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~input_o  = hps_io_hps_io_usb1_inst_D5;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~input_o  = hps_io_hps_io_usb1_inst_D6;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~input_o  = hps_io_hps_io_usb1_inst_D7;

assign \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o  = hps_io_hps_io_i2c0_inst_SDA;

assign \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o  = hps_io_hps_io_i2c0_inst_SCL;

assign \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o  = hps_io_hps_io_i2c1_inst_SDA;

assign \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o  = hps_io_hps_io_i2c1_inst_SCL;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO09;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO35;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO40;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO41;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO48;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO53;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO54;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO61;

assign \hps_f2h_irq0_irq[0]~input_o  = hps_f2h_irq0_irq[0];

assign \hps_f2h_irq0_irq[1]~input_o  = hps_f2h_irq0_irq[1];

assign \hps_f2h_irq0_irq[2]~input_o  = hps_f2h_irq0_irq[2];

assign \hps_f2h_irq0_irq[3]~input_o  = hps_f2h_irq0_irq[3];

assign \hps_f2h_irq0_irq[4]~input_o  = hps_f2h_irq0_irq[4];

assign \hps_f2h_irq0_irq[5]~input_o  = hps_f2h_irq0_irq[5];

assign \hps_f2h_irq0_irq[6]~input_o  = hps_f2h_irq0_irq[6];

assign \hps_f2h_irq0_irq[7]~input_o  = hps_f2h_irq0_irq[7];

assign \hps_f2h_irq0_irq[8]~input_o  = hps_f2h_irq0_irq[8];

assign \hps_f2h_irq0_irq[9]~input_o  = hps_f2h_irq0_irq[9];

assign \hps_f2h_irq0_irq[10]~input_o  = hps_f2h_irq0_irq[10];

assign \hps_f2h_irq0_irq[11]~input_o  = hps_f2h_irq0_irq[11];

assign \hps_f2h_irq0_irq[12]~input_o  = hps_f2h_irq0_irq[12];

assign \hps_f2h_irq0_irq[13]~input_o  = hps_f2h_irq0_irq[13];

assign \hps_f2h_irq0_irq[14]~input_o  = hps_f2h_irq0_irq[14];

assign \hps_f2h_irq0_irq[15]~input_o  = hps_f2h_irq0_irq[15];

assign \hps_f2h_irq0_irq[16]~input_o  = hps_f2h_irq0_irq[16];

assign \hps_f2h_irq0_irq[17]~input_o  = hps_f2h_irq0_irq[17];

assign \hps_f2h_irq0_irq[18]~input_o  = hps_f2h_irq0_irq[18];

assign \hps_f2h_irq0_irq[19]~input_o  = hps_f2h_irq0_irq[19];

assign \hps_f2h_irq0_irq[20]~input_o  = hps_f2h_irq0_irq[20];

assign \hps_f2h_irq0_irq[21]~input_o  = hps_f2h_irq0_irq[21];

assign \hps_f2h_irq0_irq[22]~input_o  = hps_f2h_irq0_irq[22];

assign \hps_f2h_irq0_irq[23]~input_o  = hps_f2h_irq0_irq[23];

assign \hps_f2h_irq0_irq[24]~input_o  = hps_f2h_irq0_irq[24];

assign \hps_f2h_irq0_irq[25]~input_o  = hps_f2h_irq0_irq[25];

assign \hps_f2h_irq0_irq[26]~input_o  = hps_f2h_irq0_irq[26];

assign \hps_f2h_irq0_irq[27]~input_o  = hps_f2h_irq0_irq[27];

assign \hps_f2h_irq0_irq[28]~input_o  = hps_f2h_irq0_irq[28];

assign \hps_f2h_irq0_irq[29]~input_o  = hps_f2h_irq0_irq[29];

assign \hps_f2h_irq0_irq[30]~input_o  = hps_f2h_irq0_irq[30];

assign \hps_f2h_irq0_irq[31]~input_o  = hps_f2h_irq0_irq[31];

assign \hps_io_hps_io_emac1_inst_RXD0~input_o  = hps_io_hps_io_emac1_inst_RXD0;

assign \hps_io_hps_io_emac1_inst_RXD1~input_o  = hps_io_hps_io_emac1_inst_RXD1;

assign \hps_io_hps_io_emac1_inst_RXD2~input_o  = hps_io_hps_io_emac1_inst_RXD2;

assign \hps_io_hps_io_emac1_inst_RXD3~input_o  = hps_io_hps_io_emac1_inst_RXD3;

assign \hps_io_hps_io_emac1_inst_RX_CLK~input_o  = hps_io_hps_io_emac1_inst_RX_CLK;

assign \hps_io_hps_io_emac1_inst_RX_CTL~input_o  = hps_io_hps_io_emac1_inst_RX_CTL;

assign \hps_io_hps_io_spim1_inst_MISO~input_o  = hps_io_hps_io_spim1_inst_MISO;

assign \hps_io_hps_io_uart0_inst_RX~input_o  = hps_io_hps_io_uart0_inst_RX;

assign \hps_io_hps_io_usb1_inst_CLK~input_o  = hps_io_hps_io_usb1_inst_CLK;

assign \hps_io_hps_io_usb1_inst_DIR~input_o  = hps_io_hps_io_usb1_inst_DIR;

assign \hps_io_hps_io_usb1_inst_NXT~input_o  = hps_io_hps_io_usb1_inst_NXT;

assign \memory_oct_rzqin~input_o  = memory_oct_rzqin;

assign \onchip_sram_s2_address[13]~input_o  = onchip_sram_s2_address[13];

assign \onchip_sram_s2_chipselect~input_o  = onchip_sram_s2_chipselect;

assign \onchip_sram_s2_write~input_o  = onchip_sram_s2_write;

assign \onchip_sram_clk2_clk~input_o  = onchip_sram_clk2_clk;

assign \onchip_sram_reset2_reset_req~input_o  = onchip_sram_reset2_reset_req;

assign \onchip_sram_s2_clken~input_o  = onchip_sram_s2_clken;

assign \onchip_sram_s2_writedata[0]~input_o  = onchip_sram_s2_writedata[0];

assign \onchip_sram_s2_address[0]~input_o  = onchip_sram_s2_address[0];

assign \onchip_sram_s2_address[1]~input_o  = onchip_sram_s2_address[1];

assign \onchip_sram_s2_address[2]~input_o  = onchip_sram_s2_address[2];

assign \onchip_sram_s2_address[3]~input_o  = onchip_sram_s2_address[3];

assign \onchip_sram_s2_address[4]~input_o  = onchip_sram_s2_address[4];

assign \onchip_sram_s2_address[5]~input_o  = onchip_sram_s2_address[5];

assign \onchip_sram_s2_address[6]~input_o  = onchip_sram_s2_address[6];

assign \onchip_sram_s2_address[7]~input_o  = onchip_sram_s2_address[7];

assign \onchip_sram_s2_address[8]~input_o  = onchip_sram_s2_address[8];

assign \onchip_sram_s2_address[9]~input_o  = onchip_sram_s2_address[9];

assign \onchip_sram_s2_address[10]~input_o  = onchip_sram_s2_address[10];

assign \onchip_sram_s2_address[11]~input_o  = onchip_sram_s2_address[11];

assign \onchip_sram_s2_address[12]~input_o  = onchip_sram_s2_address[12];

assign \onchip_sram_s2_byteenable[0]~input_o  = onchip_sram_s2_byteenable[0];

assign \onchip_sram_s2_writedata[1]~input_o  = onchip_sram_s2_writedata[1];

assign \onchip_sram_s2_writedata[2]~input_o  = onchip_sram_s2_writedata[2];

assign \onchip_sram_s2_writedata[3]~input_o  = onchip_sram_s2_writedata[3];

assign \onchip_sram_s2_writedata[4]~input_o  = onchip_sram_s2_writedata[4];

assign \onchip_sram_s2_writedata[5]~input_o  = onchip_sram_s2_writedata[5];

assign \onchip_sram_s2_writedata[6]~input_o  = onchip_sram_s2_writedata[6];

assign \onchip_sram_s2_writedata[7]~input_o  = onchip_sram_s2_writedata[7];

assign \onchip_sram_s2_writedata[8]~input_o  = onchip_sram_s2_writedata[8];

assign \onchip_sram_s2_byteenable[1]~input_o  = onchip_sram_s2_byteenable[1];

assign \onchip_sram_s2_writedata[9]~input_o  = onchip_sram_s2_writedata[9];

assign \onchip_sram_s2_writedata[10]~input_o  = onchip_sram_s2_writedata[10];

assign \onchip_sram_s2_writedata[11]~input_o  = onchip_sram_s2_writedata[11];

assign \onchip_sram_s2_writedata[12]~input_o  = onchip_sram_s2_writedata[12];

assign \onchip_sram_s2_writedata[13]~input_o  = onchip_sram_s2_writedata[13];

assign \onchip_sram_s2_writedata[14]~input_o  = onchip_sram_s2_writedata[14];

assign \onchip_sram_s2_writedata[15]~input_o  = onchip_sram_s2_writedata[15];

assign \onchip_sram_s2_writedata[16]~input_o  = onchip_sram_s2_writedata[16];

assign \onchip_sram_s2_byteenable[2]~input_o  = onchip_sram_s2_byteenable[2];

assign \onchip_sram_s2_writedata[17]~input_o  = onchip_sram_s2_writedata[17];

assign \onchip_sram_s2_writedata[18]~input_o  = onchip_sram_s2_writedata[18];

assign \onchip_sram_s2_writedata[19]~input_o  = onchip_sram_s2_writedata[19];

assign \onchip_sram_s2_writedata[20]~input_o  = onchip_sram_s2_writedata[20];

assign \onchip_sram_s2_writedata[21]~input_o  = onchip_sram_s2_writedata[21];

assign \onchip_sram_s2_writedata[22]~input_o  = onchip_sram_s2_writedata[22];

assign \onchip_sram_s2_writedata[23]~input_o  = onchip_sram_s2_writedata[23];

assign \onchip_sram_s2_writedata[24]~input_o  = onchip_sram_s2_writedata[24];

assign \onchip_sram_s2_byteenable[3]~input_o  = onchip_sram_s2_byteenable[3];

assign \onchip_sram_s2_writedata[25]~input_o  = onchip_sram_s2_writedata[25];

assign \onchip_sram_s2_writedata[26]~input_o  = onchip_sram_s2_writedata[26];

assign \onchip_sram_s2_writedata[27]~input_o  = onchip_sram_s2_writedata[27];

assign \onchip_sram_s2_writedata[28]~input_o  = onchip_sram_s2_writedata[28];

assign \onchip_sram_s2_writedata[29]~input_o  = onchip_sram_s2_writedata[29];

assign \onchip_sram_s2_writedata[30]~input_o  = onchip_sram_s2_writedata[30];

assign \onchip_sram_s2_writedata[31]~input_o  = onchip_sram_s2_writedata[31];

assign \system_pll_ref_clk_clk~input_o  = system_pll_ref_clk_clk;

assign \system_pll_ref_reset_reset~input_o  = system_pll_ref_reset_reset;

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck_n),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[36] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[37] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_spim1_inst_MOSI),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .shift_series_termination_control = "false";

assign hps_io_hps_io_emac1_inst_TX_CLK = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;

assign hps_io_hps_io_emac1_inst_TXD0 = \arm_a9_hps|hps_io|border|emac1_inst~emac_phy_txd ;

assign hps_io_hps_io_emac1_inst_TXD1 = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;

assign hps_io_hps_io_emac1_inst_TXD2 = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;

assign hps_io_hps_io_emac1_inst_TXD3 = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;

assign hps_io_hps_io_emac1_inst_MDC = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;

assign hps_io_hps_io_emac1_inst_TX_CTL = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;

assign hps_io_hps_io_qspi_inst_SS0 = \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;

assign hps_io_hps_io_qspi_inst_CLK = \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SCLK ;

assign hps_io_hps_io_sdio_inst_CLK = \arm_a9_hps|hps_io|border|sdio_inst~sdmmc_cclk ;

assign hps_io_hps_io_usb1_inst_STP = \arm_a9_hps|hps_io|border|usb1_inst~usb_ulpi_stp ;

assign hps_io_hps_io_spim1_inst_CLK = \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;

assign hps_io_hps_io_spim1_inst_SS0 = \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;

assign hps_io_hps_io_uart0_inst_TX = \arm_a9_hps|hps_io|border|uart0_inst~uart_txd ;

assign memory_mem_a[0] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;

assign memory_mem_a[1] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;

assign memory_mem_a[2] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;

assign memory_mem_a[3] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;

assign memory_mem_a[4] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;

assign memory_mem_a[5] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;

assign memory_mem_a[6] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;

assign memory_mem_a[7] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;

assign memory_mem_a[8] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;

assign memory_mem_a[9] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;

assign memory_mem_a[10] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;

assign memory_mem_a[11] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;

assign memory_mem_a[12] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;

assign memory_mem_a[13] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;

assign memory_mem_a[14] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;

assign memory_mem_ba[0] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;

assign memory_mem_ba[1] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;

assign memory_mem_ba[2] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;

assign memory_mem_cke = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;

assign memory_mem_cs_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;

assign memory_mem_ras_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;

assign memory_mem_cas_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;

assign memory_mem_we_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;

assign memory_mem_reset_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;

assign memory_mem_odt = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;

assign onchip_sram_s2_readdata[0] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w0_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[1] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w1_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[2] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w2_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[3] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w3_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[4] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w4_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[5] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w5_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[6] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w6_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[7] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w7_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[8] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w8_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[9] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w9_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[10] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w10_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[11] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w11_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[12] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w12_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[13] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w13_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[14] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w14_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[15] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w15_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[16] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w16_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[17] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w17_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[18] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w18_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[19] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w19_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[20] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w20_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[21] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w21_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[22] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w22_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[23] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w23_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[24] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w24_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[25] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w25_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[26] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w26_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[27] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w27_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[28] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w28_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[29] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w29_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[30] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w30_n0_mux_dataout~0_combout ;

assign onchip_sram_s2_readdata[31] = \onchip_sram|the_altsyncram|auto_generated|mux5|l1_w31_n0_mux_dataout~0_combout ;

assign sdram_clk_clk = \system_pll|sys_pll|altera_pll_i|outclk_wire[1] ;

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[0] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[1] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_emac1_inst_MDIO),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[2] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[3] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO0),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[4] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[5] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO1),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[6] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[7] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO2),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[8] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[9] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO3),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[10] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[11] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_CMD),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[12] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[13] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D0),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[14] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[15] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D1),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[16] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[17] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D2),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[18] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[19] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D3),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[20] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[21] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D0),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[22] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[23] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D1),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[24] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[25] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D2),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[26] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[27] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D3),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[28] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[29] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D4),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[30] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[31] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D5),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[32] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[33] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D6),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[34] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[35] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D7),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[38] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c0_inst_SDA),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[39] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c0_inst_SCL),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[40] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c1_inst_SDA),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[41] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c1_inst_SCL),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[42] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[43] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO09),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[44] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[45] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO35),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[46] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[47] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO40),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[48] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[49] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO41),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[50] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[51] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO48),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[52] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[53] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO53),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[54] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[55] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO54),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[56] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[57] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO61),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[4]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[5]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[6]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[7]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[8]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[9]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[10]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[11]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[12]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[13]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[14]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[15]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[16]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[17]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[18]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[19]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[20]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[21]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[22]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[23]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[24]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[25]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[26]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[27]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[28]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[29]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[30]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[31]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

assign \onchip_sram_reset2_reset~input_o  = onchip_sram_reset2_reset;

endmodule

module Computer_System_altera_reset_controller (
	h2f_rst_n_0,
	outclk_wire_0,
	locked_wire_0,
	r_early_rst1,
	r_sync_rst1)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	outclk_wire_0;
input 	locked_wire_0;
output 	r_early_rst1;
output 	r_sync_rst1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \merged_reset~0_combout ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \always2~0_combout ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;


Computer_System_altera_reset_synchronizer_2 alt_rst_req_sync_uq1(
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

Computer_System_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.merged_reset(\merged_reset~0_combout ));

cyclonev_lcell_comb \merged_reset~0 (
	.dataa(!h2f_rst_n_0),
	.datab(!locked_wire_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\merged_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_reset~0 .extended_lut = "off";
defparam \merged_reset~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \merged_reset~0 .shared_arith = "off";

dffeas r_early_rst(
	.clk(outclk_wire_0),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas r_sync_rst(
	.clk(outclk_wire_0),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(outclk_wire_0),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(outclk_wire_0),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(outclk_wire_0),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h7373737373737373;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_reset_controller_1 (
	h2f_rst_n_0,
	outclk_wire_0,
	altera_reset_synchronizer_int_chain_out)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	outclk_wire_0;
output 	altera_reset_synchronizer_int_chain_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.h2f_rst_n_0(h2f_rst_n_0),
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out));

endmodule

module Computer_System_altera_reset_synchronizer_1 (
	h2f_rst_n_0,
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_altera_reset_synchronizer_2 (
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_altera_reset_synchronizer_3 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	merged_reset)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_ARM_A9_HPS (
	h2f_rst_n_0,
	f2h_ARREADY_0,
	f2h_AWREADY_0,
	f2h_BVALID_0,
	f2h_RVALID_0,
	f2h_WREADY_0,
	f2h_RDATA_0,
	f2h_RDATA_1,
	f2h_RDATA_2,
	f2h_RDATA_3,
	f2h_RDATA_4,
	f2h_RDATA_5,
	f2h_RDATA_6,
	f2h_RDATA_7,
	f2h_RDATA_8,
	f2h_RDATA_9,
	f2h_RDATA_10,
	f2h_RDATA_11,
	f2h_RDATA_12,
	f2h_RDATA_13,
	f2h_RDATA_14,
	f2h_RDATA_15,
	f2h_RDATA_16,
	f2h_RDATA_17,
	f2h_RDATA_18,
	f2h_RDATA_19,
	f2h_RDATA_20,
	f2h_RDATA_21,
	f2h_RDATA_22,
	f2h_RDATA_23,
	f2h_RDATA_24,
	f2h_RDATA_25,
	f2h_RDATA_26,
	f2h_RDATA_27,
	f2h_RDATA_28,
	f2h_RDATA_29,
	f2h_RDATA_30,
	f2h_RDATA_31,
	f2h_RDATA_32,
	f2h_RDATA_33,
	f2h_RDATA_34,
	f2h_RDATA_35,
	f2h_RDATA_36,
	f2h_RDATA_37,
	f2h_RDATA_38,
	f2h_RDATA_39,
	f2h_RDATA_40,
	f2h_RDATA_41,
	f2h_RDATA_42,
	f2h_RDATA_43,
	f2h_RDATA_44,
	f2h_RDATA_45,
	f2h_RDATA_46,
	f2h_RDATA_47,
	f2h_RDATA_48,
	f2h_RDATA_49,
	f2h_RDATA_50,
	f2h_RDATA_51,
	f2h_RDATA_52,
	f2h_RDATA_53,
	f2h_RDATA_54,
	f2h_RDATA_55,
	f2h_RDATA_56,
	f2h_RDATA_57,
	f2h_RDATA_58,
	f2h_RDATA_59,
	f2h_RDATA_60,
	f2h_RDATA_61,
	f2h_RDATA_62,
	f2h_RDATA_63,
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	saved_grant_0,
	arvalid,
	saved_grant_1,
	awvalid,
	bready,
	wvalid,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	src_payload50,
	src_payload51,
	src_payload52,
	src_payload53,
	src_payload54,
	src_payload55,
	src_payload56,
	src_payload57,
	src_payload58,
	src_payload59,
	ShiftLeft1,
	ShiftLeft11,
	ShiftLeft12,
	ShiftLeft13,
	ShiftLeft14,
	ShiftLeft15,
	ShiftLeft16,
	ShiftLeft17,
	ShiftLeft18,
	ShiftLeft19,
	ShiftLeft110,
	ShiftLeft111,
	ShiftLeft112,
	ShiftLeft113,
	ShiftLeft114,
	ShiftLeft115,
	ShiftLeft116,
	ShiftLeft117,
	ShiftLeft118,
	ShiftLeft119,
	ShiftLeft120,
	ShiftLeft121,
	ShiftLeft122,
	ShiftLeft123,
	ShiftLeft124,
	ShiftLeft125,
	ShiftLeft126,
	ShiftLeft127,
	ShiftLeft128,
	ShiftLeft129,
	ShiftLeft130,
	ShiftLeft131,
	ShiftLeft132,
	ShiftLeft133,
	ShiftLeft134,
	ShiftLeft135,
	ShiftLeft136,
	ShiftLeft137,
	ShiftLeft138,
	ShiftLeft139,
	ShiftLeft140,
	ShiftLeft141,
	ShiftLeft142,
	ShiftLeft143,
	ShiftLeft144,
	ShiftLeft145,
	ShiftLeft146,
	ShiftLeft147,
	ShiftLeft148,
	ShiftLeft149,
	ShiftLeft150,
	ShiftLeft151,
	ShiftLeft152,
	ShiftLeft153,
	ShiftLeft154,
	ShiftLeft155,
	ShiftLeft156,
	ShiftLeft157,
	ShiftLeft158,
	ShiftLeft159,
	ShiftLeft160,
	ShiftLeft161,
	ShiftLeft162,
	ShiftLeft163,
	ShiftLeft0,
	ShiftLeft01,
	ShiftLeft02,
	ShiftLeft03,
	ShiftLeft04,
	ShiftLeft05,
	ShiftLeft06,
	ShiftLeft07,
	cmd_sink_ready,
	nonposted_cmd_accepted,
	WideOr1,
	src_payload_0,
	WideOr11,
	nonposted_cmd_accepted1,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_0,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	src_data_18,
	src_data_19,
	src_data_20,
	src_data_21,
	src_data_22,
	src_data_23,
	src_data_24,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	src_data_29,
	src_data_30,
	src_data_31,
	src_data_881,
	src_data_891,
	src_data_901,
	src_data_911,
	src_data_921,
	src_data_931,
	src_data_941,
	src_data_951,
	src_data_961,
	src_data_971,
	src_data_981,
	src_data_991,
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim1_inst,
	spim1_inst1,
	intermediate_36,
	intermediate_37,
	uart0_inst,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	intermediate_42,
	intermediate_43,
	intermediate_44,
	intermediate_46,
	intermediate_48,
	intermediate_50,
	intermediate_52,
	intermediate_54,
	intermediate_45,
	intermediate_47,
	intermediate_49,
	intermediate_51,
	intermediate_53,
	intermediate_55,
	intermediate_56,
	intermediate_57,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO35_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO41_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO53_0,
	hps_io_gpio_inst_GPIO54_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_f2h_irq0_irq_0,
	hps_f2h_irq0_irq_1,
	hps_f2h_irq0_irq_2,
	hps_f2h_irq0_irq_3,
	hps_f2h_irq0_irq_4,
	hps_f2h_irq0_irq_5,
	hps_f2h_irq0_irq_6,
	hps_f2h_irq0_irq_7,
	hps_f2h_irq0_irq_8,
	hps_f2h_irq0_irq_9,
	hps_f2h_irq0_irq_10,
	hps_f2h_irq0_irq_11,
	hps_f2h_irq0_irq_12,
	hps_f2h_irq0_irq_13,
	hps_f2h_irq0_irq_14,
	hps_f2h_irq0_irq_15,
	hps_f2h_irq0_irq_16,
	hps_f2h_irq0_irq_17,
	hps_f2h_irq0_irq_18,
	hps_f2h_irq0_irq_19,
	hps_f2h_irq0_irq_20,
	hps_f2h_irq0_irq_21,
	hps_f2h_irq0_irq_22,
	hps_f2h_irq0_irq_23,
	hps_f2h_irq0_irq_24,
	hps_f2h_irq0_irq_25,
	hps_f2h_irq0_irq_26,
	hps_f2h_irq0_irq_27,
	hps_f2h_irq0_irq_28,
	hps_f2h_irq0_irq_29,
	hps_f2h_irq0_irq_30,
	hps_f2h_irq0_irq_31,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	h2f_rst_n_0;
output 	f2h_ARREADY_0;
output 	f2h_AWREADY_0;
output 	f2h_BVALID_0;
output 	f2h_RVALID_0;
output 	f2h_WREADY_0;
output 	f2h_RDATA_0;
output 	f2h_RDATA_1;
output 	f2h_RDATA_2;
output 	f2h_RDATA_3;
output 	f2h_RDATA_4;
output 	f2h_RDATA_5;
output 	f2h_RDATA_6;
output 	f2h_RDATA_7;
output 	f2h_RDATA_8;
output 	f2h_RDATA_9;
output 	f2h_RDATA_10;
output 	f2h_RDATA_11;
output 	f2h_RDATA_12;
output 	f2h_RDATA_13;
output 	f2h_RDATA_14;
output 	f2h_RDATA_15;
output 	f2h_RDATA_16;
output 	f2h_RDATA_17;
output 	f2h_RDATA_18;
output 	f2h_RDATA_19;
output 	f2h_RDATA_20;
output 	f2h_RDATA_21;
output 	f2h_RDATA_22;
output 	f2h_RDATA_23;
output 	f2h_RDATA_24;
output 	f2h_RDATA_25;
output 	f2h_RDATA_26;
output 	f2h_RDATA_27;
output 	f2h_RDATA_28;
output 	f2h_RDATA_29;
output 	f2h_RDATA_30;
output 	f2h_RDATA_31;
output 	f2h_RDATA_32;
output 	f2h_RDATA_33;
output 	f2h_RDATA_34;
output 	f2h_RDATA_35;
output 	f2h_RDATA_36;
output 	f2h_RDATA_37;
output 	f2h_RDATA_38;
output 	f2h_RDATA_39;
output 	f2h_RDATA_40;
output 	f2h_RDATA_41;
output 	f2h_RDATA_42;
output 	f2h_RDATA_43;
output 	f2h_RDATA_44;
output 	f2h_RDATA_45;
output 	f2h_RDATA_46;
output 	f2h_RDATA_47;
output 	f2h_RDATA_48;
output 	f2h_RDATA_49;
output 	f2h_RDATA_50;
output 	f2h_RDATA_51;
output 	f2h_RDATA_52;
output 	f2h_RDATA_53;
output 	f2h_RDATA_54;
output 	f2h_RDATA_55;
output 	f2h_RDATA_56;
output 	f2h_RDATA_57;
output 	f2h_RDATA_58;
output 	f2h_RDATA_59;
output 	f2h_RDATA_60;
output 	f2h_RDATA_61;
output 	f2h_RDATA_62;
output 	f2h_RDATA_63;
output 	h2f_lw_ARVALID_0;
output 	h2f_lw_AWVALID_0;
output 	h2f_lw_BREADY_0;
output 	h2f_lw_RREADY_0;
output 	h2f_lw_WLAST_0;
output 	h2f_lw_WVALID_0;
output 	h2f_lw_ARADDR_0;
output 	h2f_lw_ARADDR_1;
output 	h2f_lw_ARADDR_2;
output 	h2f_lw_ARADDR_3;
output 	h2f_lw_ARADDR_4;
output 	h2f_lw_ARADDR_5;
output 	h2f_lw_ARBURST_0;
output 	h2f_lw_ARBURST_1;
output 	h2f_lw_ARID_0;
output 	h2f_lw_ARID_1;
output 	h2f_lw_ARID_2;
output 	h2f_lw_ARID_3;
output 	h2f_lw_ARID_4;
output 	h2f_lw_ARID_5;
output 	h2f_lw_ARID_6;
output 	h2f_lw_ARID_7;
output 	h2f_lw_ARID_8;
output 	h2f_lw_ARID_9;
output 	h2f_lw_ARID_10;
output 	h2f_lw_ARID_11;
output 	h2f_lw_ARLEN_0;
output 	h2f_lw_ARLEN_1;
output 	h2f_lw_ARLEN_2;
output 	h2f_lw_ARLEN_3;
output 	h2f_lw_ARSIZE_0;
output 	h2f_lw_ARSIZE_1;
output 	h2f_lw_ARSIZE_2;
output 	h2f_lw_AWADDR_0;
output 	h2f_lw_AWADDR_1;
output 	h2f_lw_AWADDR_2;
output 	h2f_lw_AWADDR_3;
output 	h2f_lw_AWADDR_4;
output 	h2f_lw_AWADDR_5;
output 	h2f_lw_AWBURST_0;
output 	h2f_lw_AWBURST_1;
output 	h2f_lw_AWID_0;
output 	h2f_lw_AWID_1;
output 	h2f_lw_AWID_2;
output 	h2f_lw_AWID_3;
output 	h2f_lw_AWID_4;
output 	h2f_lw_AWID_5;
output 	h2f_lw_AWID_6;
output 	h2f_lw_AWID_7;
output 	h2f_lw_AWID_8;
output 	h2f_lw_AWID_9;
output 	h2f_lw_AWID_10;
output 	h2f_lw_AWID_11;
output 	h2f_lw_AWLEN_0;
output 	h2f_lw_AWLEN_1;
output 	h2f_lw_AWLEN_2;
output 	h2f_lw_AWLEN_3;
output 	h2f_lw_AWSIZE_0;
output 	h2f_lw_AWSIZE_1;
output 	h2f_lw_AWSIZE_2;
output 	h2f_lw_WDATA_0;
output 	h2f_lw_WDATA_1;
output 	h2f_lw_WDATA_2;
output 	h2f_lw_WDATA_3;
output 	h2f_lw_WDATA_4;
output 	h2f_lw_WDATA_5;
output 	h2f_lw_WDATA_6;
output 	h2f_lw_WDATA_7;
output 	h2f_lw_WDATA_8;
output 	h2f_lw_WDATA_9;
output 	h2f_lw_WDATA_10;
output 	h2f_lw_WDATA_11;
output 	h2f_lw_WDATA_12;
output 	h2f_lw_WDATA_13;
output 	h2f_lw_WDATA_14;
output 	h2f_lw_WDATA_15;
output 	h2f_lw_WDATA_16;
output 	h2f_lw_WDATA_17;
output 	h2f_lw_WDATA_18;
output 	h2f_lw_WDATA_19;
output 	h2f_lw_WDATA_20;
output 	h2f_lw_WDATA_21;
output 	h2f_lw_WDATA_22;
output 	h2f_lw_WDATA_23;
output 	h2f_lw_WDATA_24;
output 	h2f_lw_WDATA_25;
output 	h2f_lw_WDATA_26;
output 	h2f_lw_WDATA_27;
output 	h2f_lw_WDATA_28;
output 	h2f_lw_WDATA_29;
output 	h2f_lw_WDATA_30;
output 	h2f_lw_WDATA_31;
output 	h2f_lw_WSTRB_0;
output 	h2f_lw_WSTRB_1;
output 	h2f_lw_WSTRB_2;
output 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	saved_grant_0;
input 	arvalid;
input 	saved_grant_1;
input 	awvalid;
input 	bready;
input 	wvalid;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	src_payload44;
input 	src_payload45;
input 	src_payload46;
input 	src_payload47;
input 	src_payload48;
input 	src_payload49;
input 	src_payload50;
input 	src_payload51;
input 	src_payload52;
input 	src_payload53;
input 	src_payload54;
input 	src_payload55;
input 	src_payload56;
input 	src_payload57;
input 	src_payload58;
input 	src_payload59;
input 	ShiftLeft1;
input 	ShiftLeft11;
input 	ShiftLeft12;
input 	ShiftLeft13;
input 	ShiftLeft14;
input 	ShiftLeft15;
input 	ShiftLeft16;
input 	ShiftLeft17;
input 	ShiftLeft18;
input 	ShiftLeft19;
input 	ShiftLeft110;
input 	ShiftLeft111;
input 	ShiftLeft112;
input 	ShiftLeft113;
input 	ShiftLeft114;
input 	ShiftLeft115;
input 	ShiftLeft116;
input 	ShiftLeft117;
input 	ShiftLeft118;
input 	ShiftLeft119;
input 	ShiftLeft120;
input 	ShiftLeft121;
input 	ShiftLeft122;
input 	ShiftLeft123;
input 	ShiftLeft124;
input 	ShiftLeft125;
input 	ShiftLeft126;
input 	ShiftLeft127;
input 	ShiftLeft128;
input 	ShiftLeft129;
input 	ShiftLeft130;
input 	ShiftLeft131;
input 	ShiftLeft132;
input 	ShiftLeft133;
input 	ShiftLeft134;
input 	ShiftLeft135;
input 	ShiftLeft136;
input 	ShiftLeft137;
input 	ShiftLeft138;
input 	ShiftLeft139;
input 	ShiftLeft140;
input 	ShiftLeft141;
input 	ShiftLeft142;
input 	ShiftLeft143;
input 	ShiftLeft144;
input 	ShiftLeft145;
input 	ShiftLeft146;
input 	ShiftLeft147;
input 	ShiftLeft148;
input 	ShiftLeft149;
input 	ShiftLeft150;
input 	ShiftLeft151;
input 	ShiftLeft152;
input 	ShiftLeft153;
input 	ShiftLeft154;
input 	ShiftLeft155;
input 	ShiftLeft156;
input 	ShiftLeft157;
input 	ShiftLeft158;
input 	ShiftLeft159;
input 	ShiftLeft160;
input 	ShiftLeft161;
input 	ShiftLeft162;
input 	ShiftLeft163;
input 	ShiftLeft0;
input 	ShiftLeft01;
input 	ShiftLeft02;
input 	ShiftLeft03;
input 	ShiftLeft04;
input 	ShiftLeft05;
input 	ShiftLeft06;
input 	ShiftLeft07;
input 	cmd_sink_ready;
input 	nonposted_cmd_accepted;
input 	WideOr1;
input 	src_payload_0;
input 	WideOr11;
input 	nonposted_cmd_accepted1;
input 	src_data_88;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_0;
input 	src_data_1;
input 	src_data_2;
input 	src_data_3;
input 	src_data_4;
input 	src_data_5;
input 	src_data_6;
input 	src_data_7;
input 	src_data_8;
input 	src_data_9;
input 	src_data_10;
input 	src_data_11;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_data_17;
input 	src_data_18;
input 	src_data_19;
input 	src_data_20;
input 	src_data_21;
input 	src_data_22;
input 	src_data_23;
input 	src_data_24;
input 	src_data_25;
input 	src_data_26;
input 	src_data_27;
input 	src_data_28;
input 	src_data_29;
input 	src_data_30;
input 	src_data_31;
input 	src_data_881;
input 	src_data_891;
input 	src_data_901;
input 	src_data_911;
input 	src_data_921;
input 	src_data_931;
input 	src_data_941;
input 	src_data_951;
input 	src_data_961;
input 	src_data_971;
input 	src_data_981;
input 	src_data_991;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	uart0_inst;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	intermediate_42;
output 	intermediate_43;
output 	intermediate_44;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_50;
output 	intermediate_52;
output 	intermediate_54;
output 	intermediate_45;
output 	intermediate_47;
output 	intermediate_49;
output 	intermediate_51;
output 	intermediate_53;
output 	intermediate_55;
output 	intermediate_56;
output 	intermediate_57;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO35_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO41_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO53_0;
input 	hps_io_gpio_inst_GPIO54_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_f2h_irq0_irq_0;
input 	hps_f2h_irq0_irq_1;
input 	hps_f2h_irq0_irq_2;
input 	hps_f2h_irq0_irq_3;
input 	hps_f2h_irq0_irq_4;
input 	hps_f2h_irq0_irq_5;
input 	hps_f2h_irq0_irq_6;
input 	hps_f2h_irq0_irq_7;
input 	hps_f2h_irq0_irq_8;
input 	hps_f2h_irq0_irq_9;
input 	hps_f2h_irq0_irq_10;
input 	hps_f2h_irq0_irq_11;
input 	hps_f2h_irq0_irq_12;
input 	hps_f2h_irq0_irq_13;
input 	hps_f2h_irq0_irq_14;
input 	hps_f2h_irq0_irq_15;
input 	hps_f2h_irq0_irq_16;
input 	hps_f2h_irq0_irq_17;
input 	hps_f2h_irq0_irq_18;
input 	hps_f2h_irq0_irq_19;
input 	hps_f2h_irq0_irq_20;
input 	hps_f2h_irq0_irq_21;
input 	hps_f2h_irq0_irq_22;
input 	hps_f2h_irq0_irq_23;
input 	hps_f2h_irq0_irq_24;
input 	hps_f2h_irq0_irq_25;
input 	hps_f2h_irq0_irq_26;
input 	hps_f2h_irq0_irq_27;
input 	hps_f2h_irq0_irq_28;
input 	hps_f2h_irq0_irq_29;
input 	hps_f2h_irq0_irq_30;
input 	hps_f2h_irq0_irq_31;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_ARM_A9_HPS_hps_io hps_io(
	.emac1_inst(emac1_inst),
	.emac1_inst1(emac1_inst1),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.emac1_inst2(emac1_inst2),
	.emac1_inst3(emac1_inst3),
	.emac1_inst4(emac1_inst4),
	.emac1_inst5(emac1_inst5),
	.emac1_inst6(emac1_inst6),
	.qspi_inst(qspi_inst),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.qspi_inst1(qspi_inst1),
	.sdio_inst(sdio_inst),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.usb1_inst(usb1_inst),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.spim1_inst(spim1_inst),
	.spim1_inst1(spim1_inst1),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.uart0_inst(uart0_inst),
	.intermediate_39(intermediate_39),
	.intermediate_38(intermediate_38),
	.intermediate_41(intermediate_41),
	.intermediate_40(intermediate_40),
	.intermediate_42(intermediate_42),
	.intermediate_43(intermediate_43),
	.intermediate_44(intermediate_44),
	.intermediate_46(intermediate_46),
	.intermediate_48(intermediate_48),
	.intermediate_50(intermediate_50),
	.intermediate_52(intermediate_52),
	.intermediate_54(intermediate_54),
	.intermediate_45(intermediate_45),
	.intermediate_47(intermediate_47),
	.intermediate_49(intermediate_49),
	.intermediate_51(intermediate_51),
	.intermediate_53(intermediate_53),
	.intermediate_55(intermediate_55),
	.intermediate_56(intermediate_56),
	.intermediate_57(intermediate_57),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_i2c0_inst_SDA_0(hps_io_i2c0_inst_SDA_0),
	.hps_io_i2c0_inst_SCL_0(hps_io_i2c0_inst_SCL_0),
	.hps_io_i2c1_inst_SDA_0(hps_io_i2c1_inst_SDA_0),
	.hps_io_i2c1_inst_SCL_0(hps_io_i2c1_inst_SCL_0),
	.hps_io_gpio_inst_GPIO09_0(hps_io_gpio_inst_GPIO09_0),
	.hps_io_gpio_inst_GPIO35_0(hps_io_gpio_inst_GPIO35_0),
	.hps_io_gpio_inst_GPIO40_0(hps_io_gpio_inst_GPIO40_0),
	.hps_io_gpio_inst_GPIO41_0(hps_io_gpio_inst_GPIO41_0),
	.hps_io_gpio_inst_GPIO48_0(hps_io_gpio_inst_GPIO48_0),
	.hps_io_gpio_inst_GPIO53_0(hps_io_gpio_inst_GPIO53_0),
	.hps_io_gpio_inst_GPIO54_0(hps_io_gpio_inst_GPIO54_0),
	.hps_io_gpio_inst_GPIO61_0(hps_io_gpio_inst_GPIO61_0),
	.hps_io_hps_io_emac1_inst_RXD0(hps_io_hps_io_emac1_inst_RXD0),
	.hps_io_hps_io_emac1_inst_RXD1(hps_io_hps_io_emac1_inst_RXD1),
	.hps_io_hps_io_emac1_inst_RXD2(hps_io_hps_io_emac1_inst_RXD2),
	.hps_io_hps_io_emac1_inst_RXD3(hps_io_hps_io_emac1_inst_RXD3),
	.hps_io_hps_io_emac1_inst_RX_CLK(hps_io_hps_io_emac1_inst_RX_CLK),
	.hps_io_hps_io_emac1_inst_RX_CTL(hps_io_hps_io_emac1_inst_RX_CTL),
	.hps_io_hps_io_spim1_inst_MISO(hps_io_hps_io_spim1_inst_MISO),
	.hps_io_hps_io_uart0_inst_RX(hps_io_hps_io_uart0_inst_RX),
	.hps_io_hps_io_usb1_inst_CLK(hps_io_hps_io_usb1_inst_CLK),
	.hps_io_hps_io_usb1_inst_DIR(hps_io_hps_io_usb1_inst_DIR),
	.hps_io_hps_io_usb1_inst_NXT(hps_io_hps_io_usb1_inst_NXT),
	.memory_oct_rzqin(memory_oct_rzqin));

Computer_System_Computer_System_ARM_A9_HPS_fpga_interfaces fpga_interfaces(
	.h2f_rst_n({h2f_rst_n_0}),
	.f2h_ARREADY({f2h_ARREADY_0}),
	.f2h_AWREADY({f2h_AWREADY_0}),
	.f2h_BVALID({f2h_BVALID_0}),
	.f2h_RVALID({f2h_RVALID_0}),
	.f2h_WREADY({f2h_WREADY_0}),
	.f2h_RDATA({f2h_RDATA_63,f2h_RDATA_62,f2h_RDATA_61,f2h_RDATA_60,f2h_RDATA_59,f2h_RDATA_58,f2h_RDATA_57,f2h_RDATA_56,f2h_RDATA_55,f2h_RDATA_54,f2h_RDATA_53,f2h_RDATA_52,f2h_RDATA_51,f2h_RDATA_50,f2h_RDATA_49,f2h_RDATA_48,f2h_RDATA_47,f2h_RDATA_46,f2h_RDATA_45,f2h_RDATA_44,f2h_RDATA_43,
f2h_RDATA_42,f2h_RDATA_41,f2h_RDATA_40,f2h_RDATA_39,f2h_RDATA_38,f2h_RDATA_37,f2h_RDATA_36,f2h_RDATA_35,f2h_RDATA_34,f2h_RDATA_33,f2h_RDATA_32,f2h_RDATA_31,f2h_RDATA_30,f2h_RDATA_29,f2h_RDATA_28,f2h_RDATA_27,f2h_RDATA_26,f2h_RDATA_25,f2h_RDATA_24,f2h_RDATA_23,f2h_RDATA_22,
f2h_RDATA_21,f2h_RDATA_20,f2h_RDATA_19,f2h_RDATA_18,f2h_RDATA_17,f2h_RDATA_16,f2h_RDATA_15,f2h_RDATA_14,f2h_RDATA_13,f2h_RDATA_12,f2h_RDATA_11,f2h_RDATA_10,f2h_RDATA_9,f2h_RDATA_8,f2h_RDATA_7,f2h_RDATA_6,f2h_RDATA_5,f2h_RDATA_4,f2h_RDATA_3,f2h_RDATA_2,f2h_RDATA_1,f2h_RDATA_0}),
	.h2f_lw_ARVALID({h2f_lw_ARVALID_0}),
	.h2f_lw_AWVALID({h2f_lw_AWVALID_0}),
	.h2f_lw_BREADY({h2f_lw_BREADY_0}),
	.h2f_lw_RREADY({h2f_lw_RREADY_0}),
	.h2f_lw_WLAST({h2f_lw_WLAST_0}),
	.h2f_lw_WVALID({h2f_lw_WVALID_0}),
	.h2f_lw_ARADDR({h2f_lw_ARADDR_unconnected_wire_20,h2f_lw_ARADDR_unconnected_wire_19,h2f_lw_ARADDR_unconnected_wire_18,h2f_lw_ARADDR_unconnected_wire_17,h2f_lw_ARADDR_unconnected_wire_16,h2f_lw_ARADDR_unconnected_wire_15,h2f_lw_ARADDR_unconnected_wire_14,
h2f_lw_ARADDR_unconnected_wire_13,h2f_lw_ARADDR_unconnected_wire_12,h2f_lw_ARADDR_unconnected_wire_11,h2f_lw_ARADDR_unconnected_wire_10,h2f_lw_ARADDR_unconnected_wire_9,h2f_lw_ARADDR_unconnected_wire_8,h2f_lw_ARADDR_unconnected_wire_7,
h2f_lw_ARADDR_unconnected_wire_6,h2f_lw_ARADDR_5,h2f_lw_ARADDR_4,h2f_lw_ARADDR_3,h2f_lw_ARADDR_2,h2f_lw_ARADDR_1,h2f_lw_ARADDR_0}),
	.h2f_lw_ARBURST({h2f_lw_ARBURST_1,h2f_lw_ARBURST_0}),
	.h2f_lw_ARID({h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0}),
	.h2f_lw_ARLEN({h2f_lw_ARLEN_3,h2f_lw_ARLEN_2,h2f_lw_ARLEN_1,h2f_lw_ARLEN_0}),
	.h2f_lw_ARSIZE({h2f_lw_ARSIZE_2,h2f_lw_ARSIZE_1,h2f_lw_ARSIZE_0}),
	.h2f_lw_AWADDR({h2f_lw_AWADDR_unconnected_wire_20,h2f_lw_AWADDR_unconnected_wire_19,h2f_lw_AWADDR_unconnected_wire_18,h2f_lw_AWADDR_unconnected_wire_17,h2f_lw_AWADDR_unconnected_wire_16,h2f_lw_AWADDR_unconnected_wire_15,h2f_lw_AWADDR_unconnected_wire_14,
h2f_lw_AWADDR_unconnected_wire_13,h2f_lw_AWADDR_unconnected_wire_12,h2f_lw_AWADDR_unconnected_wire_11,h2f_lw_AWADDR_unconnected_wire_10,h2f_lw_AWADDR_unconnected_wire_9,h2f_lw_AWADDR_unconnected_wire_8,h2f_lw_AWADDR_unconnected_wire_7,
h2f_lw_AWADDR_unconnected_wire_6,h2f_lw_AWADDR_5,h2f_lw_AWADDR_4,h2f_lw_AWADDR_3,h2f_lw_AWADDR_2,h2f_lw_AWADDR_1,h2f_lw_AWADDR_0}),
	.h2f_lw_AWBURST({h2f_lw_AWBURST_1,h2f_lw_AWBURST_0}),
	.h2f_lw_AWID({h2f_lw_AWID_11,h2f_lw_AWID_10,h2f_lw_AWID_9,h2f_lw_AWID_8,h2f_lw_AWID_7,h2f_lw_AWID_6,h2f_lw_AWID_5,h2f_lw_AWID_4,h2f_lw_AWID_3,h2f_lw_AWID_2,h2f_lw_AWID_1,h2f_lw_AWID_0}),
	.h2f_lw_AWLEN({h2f_lw_AWLEN_3,h2f_lw_AWLEN_2,h2f_lw_AWLEN_1,h2f_lw_AWLEN_0}),
	.h2f_lw_AWSIZE({h2f_lw_AWSIZE_2,h2f_lw_AWSIZE_1,h2f_lw_AWSIZE_0}),
	.h2f_lw_WDATA({h2f_lw_WDATA_31,h2f_lw_WDATA_30,h2f_lw_WDATA_29,h2f_lw_WDATA_28,h2f_lw_WDATA_27,h2f_lw_WDATA_26,h2f_lw_WDATA_25,h2f_lw_WDATA_24,h2f_lw_WDATA_23,h2f_lw_WDATA_22,h2f_lw_WDATA_21,h2f_lw_WDATA_20,h2f_lw_WDATA_19,h2f_lw_WDATA_18,h2f_lw_WDATA_17,h2f_lw_WDATA_16,h2f_lw_WDATA_15,
h2f_lw_WDATA_14,h2f_lw_WDATA_13,h2f_lw_WDATA_12,h2f_lw_WDATA_11,h2f_lw_WDATA_10,h2f_lw_WDATA_9,h2f_lw_WDATA_8,h2f_lw_WDATA_7,h2f_lw_WDATA_6,h2f_lw_WDATA_5,h2f_lw_WDATA_4,h2f_lw_WDATA_3,h2f_lw_WDATA_2,h2f_lw_WDATA_1,h2f_lw_WDATA_0}),
	.h2f_lw_WSTRB({h2f_lw_WSTRB_3,h2f_lw_WSTRB_2,h2f_lw_WSTRB_1,h2f_lw_WSTRB_0}),
	.h2f_lw_axi_clk({outclk_wire_0}),
	.f2h_axi_clk({outclk_wire_0}),
	.h2f_axi_clk({outclk_wire_0}),
	.f2h_ARSIZE({gnd,saved_grant_0,gnd}),
	.f2h_ARPROT({gnd,saved_grant_0,gnd}),
	.f2h_ARBURST({gnd,saved_grant_0}),
	.f2h_ARVALID({arvalid}),
	.f2h_AWSIZE({gnd,saved_grant_1,gnd}),
	.f2h_AWPROT({gnd,saved_grant_1,gnd}),
	.f2h_AWLEN({saved_grant_1,saved_grant_1,saved_grant_1,saved_grant_1}),
	.f2h_AWBURST({gnd,saved_grant_1}),
	.f2h_WLAST({saved_grant_1}),
	.f2h_AWVALID({awvalid}),
	.f2h_BREADY({bready}),
	.f2h_WVALID({wvalid}),
	.f2h_ARADDR({src_payload29,src_payload28,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,
src_payload10,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload,gnd,gnd}),
	.f2h_AWADDR({src_payload59,src_payload58,src_payload57,src_payload56,src_payload55,src_payload54,src_payload53,src_payload52,src_payload51,src_payload50,src_payload49,src_payload48,src_payload47,src_payload46,src_payload45,src_payload44,src_payload43,src_payload42,src_payload41,
src_payload40,src_payload39,src_payload38,src_payload37,src_payload36,src_payload35,src_payload34,src_payload33,src_payload32,src_payload31,src_payload30,gnd,gnd}),
	.f2h_WDATA({ShiftLeft163,ShiftLeft162,ShiftLeft161,ShiftLeft160,ShiftLeft159,ShiftLeft158,ShiftLeft157,ShiftLeft156,ShiftLeft155,ShiftLeft154,ShiftLeft153,ShiftLeft152,ShiftLeft151,ShiftLeft150,ShiftLeft149,ShiftLeft148,ShiftLeft147,ShiftLeft146,ShiftLeft145,ShiftLeft144,ShiftLeft143,
ShiftLeft142,ShiftLeft141,ShiftLeft140,ShiftLeft139,ShiftLeft138,ShiftLeft137,ShiftLeft136,ShiftLeft135,ShiftLeft134,ShiftLeft133,ShiftLeft132,ShiftLeft131,ShiftLeft130,ShiftLeft129,ShiftLeft128,ShiftLeft127,ShiftLeft126,ShiftLeft125,ShiftLeft124,ShiftLeft123,ShiftLeft122,
ShiftLeft121,ShiftLeft120,ShiftLeft119,ShiftLeft118,ShiftLeft117,ShiftLeft116,ShiftLeft115,ShiftLeft114,ShiftLeft113,ShiftLeft112,ShiftLeft111,ShiftLeft110,ShiftLeft19,ShiftLeft18,ShiftLeft17,ShiftLeft16,ShiftLeft15,ShiftLeft14,ShiftLeft13,ShiftLeft12,ShiftLeft11,ShiftLeft1}),
	.f2h_WSTRB({ShiftLeft07,ShiftLeft06,ShiftLeft05,ShiftLeft04,ShiftLeft03,ShiftLeft02,ShiftLeft01,ShiftLeft0}),
	.h2f_lw_ARREADY({cmd_sink_ready}),
	.h2f_lw_AWREADY({nonposted_cmd_accepted}),
	.h2f_lw_BVALID({WideOr1}),
	.h2f_lw_RLAST({src_payload_0}),
	.h2f_lw_RVALID({WideOr11}),
	.h2f_lw_WREADY({nonposted_cmd_accepted1}),
	.h2f_lw_BID({src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,src_data_91,src_data_90,src_data_89,src_data_88}),
	.h2f_lw_RDATA({src_data_31,src_data_30,src_data_29,src_data_28,src_data_27,src_data_26,src_data_25,src_data_24,src_data_23,src_data_22,src_data_21,src_data_20,src_data_19,src_data_18,src_data_17,src_data_16,src_data_15,src_data_14,src_data_13,src_data_12,src_data_11,src_data_10,src_data_9,
src_data_8,src_data_7,src_data_6,src_data_5,src_data_4,src_data_3,src_data_2,src_data_1,src_data_0}),
	.h2f_lw_RID({src_data_991,src_data_981,src_data_971,src_data_961,src_data_951,src_data_941,src_data_931,src_data_921,src_data_911,src_data_901,src_data_891,src_data_881}),
	.f2h_irq_p0({hps_f2h_irq0_irq_31,hps_f2h_irq0_irq_30,hps_f2h_irq0_irq_29,hps_f2h_irq0_irq_28,hps_f2h_irq0_irq_27,hps_f2h_irq0_irq_26,hps_f2h_irq0_irq_25,hps_f2h_irq0_irq_24,hps_f2h_irq0_irq_23,hps_f2h_irq0_irq_22,hps_f2h_irq0_irq_21,hps_f2h_irq0_irq_20,hps_f2h_irq0_irq_19,
hps_f2h_irq0_irq_18,hps_f2h_irq0_irq_17,hps_f2h_irq0_irq_16,hps_f2h_irq0_irq_15,hps_f2h_irq0_irq_14,hps_f2h_irq0_irq_13,hps_f2h_irq0_irq_12,hps_f2h_irq0_irq_11,hps_f2h_irq0_irq_10,hps_f2h_irq0_irq_9,hps_f2h_irq0_irq_8,hps_f2h_irq0_irq_7,hps_f2h_irq0_irq_6,
hps_f2h_irq0_irq_5,hps_f2h_irq0_irq_4,hps_f2h_irq0_irq_3,hps_f2h_irq0_irq_2,hps_f2h_irq0_irq_1,hps_f2h_irq0_irq_0}));

endmodule

module Computer_System_Computer_System_ARM_A9_HPS_fpga_interfaces (
	h2f_rst_n,
	f2h_ARREADY,
	f2h_AWREADY,
	f2h_BVALID,
	f2h_RVALID,
	f2h_WREADY,
	f2h_RDATA,
	h2f_lw_ARVALID,
	h2f_lw_AWVALID,
	h2f_lw_BREADY,
	h2f_lw_RREADY,
	h2f_lw_WLAST,
	h2f_lw_WVALID,
	h2f_lw_ARADDR,
	h2f_lw_ARBURST,
	h2f_lw_ARID,
	h2f_lw_ARLEN,
	h2f_lw_ARSIZE,
	h2f_lw_AWADDR,
	h2f_lw_AWBURST,
	h2f_lw_AWID,
	h2f_lw_AWLEN,
	h2f_lw_AWSIZE,
	h2f_lw_WDATA,
	h2f_lw_WSTRB,
	h2f_lw_axi_clk,
	f2h_axi_clk,
	h2f_axi_clk,
	f2h_ARSIZE,
	f2h_ARPROT,
	f2h_ARBURST,
	f2h_ARVALID,
	f2h_AWSIZE,
	f2h_AWPROT,
	f2h_AWLEN,
	f2h_AWBURST,
	f2h_WLAST,
	f2h_AWVALID,
	f2h_BREADY,
	f2h_WVALID,
	f2h_ARADDR,
	f2h_AWADDR,
	f2h_WDATA,
	f2h_WSTRB,
	h2f_lw_ARREADY,
	h2f_lw_AWREADY,
	h2f_lw_BVALID,
	h2f_lw_RLAST,
	h2f_lw_RVALID,
	h2f_lw_WREADY,
	h2f_lw_BID,
	h2f_lw_RDATA,
	h2f_lw_RID,
	f2h_irq_p0)/* synthesis synthesis_greybox=0 */;
output 	[0:0] h2f_rst_n;
output 	[0:0] f2h_ARREADY;
output 	[0:0] f2h_AWREADY;
output 	[0:0] f2h_BVALID;
output 	[0:0] f2h_RVALID;
output 	[0:0] f2h_WREADY;
output 	[63:0] f2h_RDATA;
output 	[0:0] h2f_lw_ARVALID;
output 	[0:0] h2f_lw_AWVALID;
output 	[0:0] h2f_lw_BREADY;
output 	[0:0] h2f_lw_RREADY;
output 	[0:0] h2f_lw_WLAST;
output 	[0:0] h2f_lw_WVALID;
output 	[20:0] h2f_lw_ARADDR;
output 	[1:0] h2f_lw_ARBURST;
output 	[11:0] h2f_lw_ARID;
output 	[3:0] h2f_lw_ARLEN;
output 	[2:0] h2f_lw_ARSIZE;
output 	[20:0] h2f_lw_AWADDR;
output 	[1:0] h2f_lw_AWBURST;
output 	[11:0] h2f_lw_AWID;
output 	[3:0] h2f_lw_AWLEN;
output 	[2:0] h2f_lw_AWSIZE;
output 	[31:0] h2f_lw_WDATA;
output 	[3:0] h2f_lw_WSTRB;
input 	[0:0] h2f_lw_axi_clk;
input 	[0:0] f2h_axi_clk;
input 	[0:0] h2f_axi_clk;
input 	[2:0] f2h_ARSIZE;
input 	[2:0] f2h_ARPROT;
input 	[1:0] f2h_ARBURST;
input 	[0:0] f2h_ARVALID;
input 	[2:0] f2h_AWSIZE;
input 	[2:0] f2h_AWPROT;
input 	[3:0] f2h_AWLEN;
input 	[1:0] f2h_AWBURST;
input 	[0:0] f2h_WLAST;
input 	[0:0] f2h_AWVALID;
input 	[0:0] f2h_BREADY;
input 	[0:0] f2h_WVALID;
input 	[31:0] f2h_ARADDR;
input 	[31:0] f2h_AWADDR;
input 	[63:0] f2h_WDATA;
input 	[7:0] f2h_WSTRB;
input 	[0:0] h2f_lw_ARREADY;
input 	[0:0] h2f_lw_AWREADY;
input 	[0:0] h2f_lw_BVALID;
input 	[0:0] h2f_lw_RLAST;
input 	[0:0] h2f_lw_RVALID;
input 	[0:0] h2f_lw_WREADY;
input 	[11:0] h2f_lw_BID;
input 	[31:0] h2f_lw_RDATA;
input 	[11:0] h2f_lw_RID;
input 	[31:0] f2h_irq_p0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \debug_apb~O_P_ADDR_31 ;
wire \tpiu~trace_data ;
wire \tpiu~O_TRACE_DATA1 ;
wire \tpiu~O_TRACE_DATA2 ;
wire \tpiu~O_TRACE_DATA3 ;
wire \tpiu~O_TRACE_DATA4 ;
wire \tpiu~O_TRACE_DATA5 ;
wire \tpiu~O_TRACE_DATA6 ;
wire \tpiu~O_TRACE_DATA7 ;
wire \tpiu~O_TRACE_DATA8 ;
wire \tpiu~O_TRACE_DATA9 ;
wire \tpiu~O_TRACE_DATA10 ;
wire \tpiu~O_TRACE_DATA11 ;
wire \tpiu~O_TRACE_DATA12 ;
wire \tpiu~O_TRACE_DATA13 ;
wire \tpiu~O_TRACE_DATA14 ;
wire \tpiu~O_TRACE_DATA15 ;
wire \tpiu~O_TRACE_DATA16 ;
wire \tpiu~O_TRACE_DATA17 ;
wire \tpiu~O_TRACE_DATA18 ;
wire \tpiu~O_TRACE_DATA19 ;
wire \tpiu~O_TRACE_DATA20 ;
wire \tpiu~O_TRACE_DATA21 ;
wire \tpiu~O_TRACE_DATA22 ;
wire \tpiu~O_TRACE_DATA23 ;
wire \tpiu~O_TRACE_DATA24 ;
wire \tpiu~O_TRACE_DATA25 ;
wire \tpiu~O_TRACE_DATA26 ;
wire \tpiu~O_TRACE_DATA27 ;
wire \tpiu~O_TRACE_DATA28 ;
wire \tpiu~O_TRACE_DATA29 ;
wire \tpiu~O_TRACE_DATA30 ;
wire \tpiu~O_TRACE_DATA31 ;
wire \boot_from_fpga~fake_dout ;
wire \h2f_ARADDR[0] ;
wire \h2f_ARADDR[1] ;
wire \h2f_ARADDR[2] ;
wire \h2f_ARADDR[3] ;
wire \h2f_ARADDR[4] ;
wire \h2f_ARADDR[5] ;
wire \h2f_ARADDR[6] ;
wire \h2f_ARADDR[7] ;
wire \h2f_ARADDR[8] ;
wire \h2f_ARADDR[9] ;
wire \h2f_ARADDR[10] ;
wire \h2f_ARADDR[11] ;
wire \h2f_ARADDR[12] ;
wire \h2f_ARADDR[13] ;
wire \h2f_ARADDR[14] ;
wire \h2f_ARADDR[15] ;
wire \h2f_ARADDR[16] ;
wire \h2f_ARADDR[17] ;
wire \h2f_ARADDR[18] ;
wire \h2f_ARADDR[19] ;
wire \h2f_ARADDR[20] ;
wire \h2f_ARADDR[21] ;
wire \h2f_ARADDR[22] ;
wire \h2f_ARADDR[23] ;
wire \h2f_ARADDR[24] ;
wire \h2f_ARADDR[25] ;
wire \h2f_ARADDR[26] ;
wire \h2f_ARADDR[27] ;
wire \h2f_ARADDR[28] ;
wire \h2f_ARADDR[29] ;
wire \f2sdram~O_BONDING_OUT_10 ;
wire \f2sdram~O_BONDING_OUT_11 ;
wire \f2sdram~O_BONDING_OUT_12 ;
wire \f2sdram~O_BONDING_OUT_13 ;
wire \interrupts~fake_dout ;
wire \clocks_resets~h2f_cold_rst_n ;
wire \h2f_lw_ARADDR[6] ;
wire \h2f_lw_ARADDR[7] ;
wire \h2f_lw_ARADDR[8] ;
wire \h2f_lw_ARADDR[9] ;
wire \h2f_lw_ARADDR[10] ;
wire \h2f_lw_ARADDR[11] ;
wire \h2f_lw_ARADDR[12] ;
wire \h2f_lw_ARADDR[13] ;
wire \h2f_lw_ARADDR[14] ;
wire \h2f_lw_ARADDR[15] ;
wire \h2f_lw_ARADDR[16] ;
wire \h2f_lw_ARADDR[17] ;
wire \h2f_lw_ARADDR[18] ;
wire \h2f_lw_ARADDR[19] ;
wire \h2f_lw_ARADDR[20] ;

wire [31:0] tpiu_TRACE_DATA_bus;
wire [29:0] hps2fpga_ARADDR_bus;
wire [3:0] f2sdram_BONDING_OUT_1_bus;
wire [127:0] fpga2hps_RDATA_bus;
wire [20:0] hps2fpga_light_weight_ARADDR_bus;
wire [1:0] hps2fpga_light_weight_ARBURST_bus;
wire [11:0] hps2fpga_light_weight_ARID_bus;
wire [3:0] hps2fpga_light_weight_ARLEN_bus;
wire [2:0] hps2fpga_light_weight_ARSIZE_bus;
wire [20:0] hps2fpga_light_weight_AWADDR_bus;
wire [1:0] hps2fpga_light_weight_AWBURST_bus;
wire [11:0] hps2fpga_light_weight_AWID_bus;
wire [3:0] hps2fpga_light_weight_AWLEN_bus;
wire [2:0] hps2fpga_light_weight_AWSIZE_bus;
wire [31:0] hps2fpga_light_weight_WDATA_bus;
wire [3:0] hps2fpga_light_weight_WSTRB_bus;

assign \tpiu~trace_data  = tpiu_TRACE_DATA_bus[0];
assign \tpiu~O_TRACE_DATA1  = tpiu_TRACE_DATA_bus[1];
assign \tpiu~O_TRACE_DATA2  = tpiu_TRACE_DATA_bus[2];
assign \tpiu~O_TRACE_DATA3  = tpiu_TRACE_DATA_bus[3];
assign \tpiu~O_TRACE_DATA4  = tpiu_TRACE_DATA_bus[4];
assign \tpiu~O_TRACE_DATA5  = tpiu_TRACE_DATA_bus[5];
assign \tpiu~O_TRACE_DATA6  = tpiu_TRACE_DATA_bus[6];
assign \tpiu~O_TRACE_DATA7  = tpiu_TRACE_DATA_bus[7];
assign \tpiu~O_TRACE_DATA8  = tpiu_TRACE_DATA_bus[8];
assign \tpiu~O_TRACE_DATA9  = tpiu_TRACE_DATA_bus[9];
assign \tpiu~O_TRACE_DATA10  = tpiu_TRACE_DATA_bus[10];
assign \tpiu~O_TRACE_DATA11  = tpiu_TRACE_DATA_bus[11];
assign \tpiu~O_TRACE_DATA12  = tpiu_TRACE_DATA_bus[12];
assign \tpiu~O_TRACE_DATA13  = tpiu_TRACE_DATA_bus[13];
assign \tpiu~O_TRACE_DATA14  = tpiu_TRACE_DATA_bus[14];
assign \tpiu~O_TRACE_DATA15  = tpiu_TRACE_DATA_bus[15];
assign \tpiu~O_TRACE_DATA16  = tpiu_TRACE_DATA_bus[16];
assign \tpiu~O_TRACE_DATA17  = tpiu_TRACE_DATA_bus[17];
assign \tpiu~O_TRACE_DATA18  = tpiu_TRACE_DATA_bus[18];
assign \tpiu~O_TRACE_DATA19  = tpiu_TRACE_DATA_bus[19];
assign \tpiu~O_TRACE_DATA20  = tpiu_TRACE_DATA_bus[20];
assign \tpiu~O_TRACE_DATA21  = tpiu_TRACE_DATA_bus[21];
assign \tpiu~O_TRACE_DATA22  = tpiu_TRACE_DATA_bus[22];
assign \tpiu~O_TRACE_DATA23  = tpiu_TRACE_DATA_bus[23];
assign \tpiu~O_TRACE_DATA24  = tpiu_TRACE_DATA_bus[24];
assign \tpiu~O_TRACE_DATA25  = tpiu_TRACE_DATA_bus[25];
assign \tpiu~O_TRACE_DATA26  = tpiu_TRACE_DATA_bus[26];
assign \tpiu~O_TRACE_DATA27  = tpiu_TRACE_DATA_bus[27];
assign \tpiu~O_TRACE_DATA28  = tpiu_TRACE_DATA_bus[28];
assign \tpiu~O_TRACE_DATA29  = tpiu_TRACE_DATA_bus[29];
assign \tpiu~O_TRACE_DATA30  = tpiu_TRACE_DATA_bus[30];
assign \tpiu~O_TRACE_DATA31  = tpiu_TRACE_DATA_bus[31];

assign \h2f_ARADDR[0]  = hps2fpga_ARADDR_bus[0];
assign \h2f_ARADDR[1]  = hps2fpga_ARADDR_bus[1];
assign \h2f_ARADDR[2]  = hps2fpga_ARADDR_bus[2];
assign \h2f_ARADDR[3]  = hps2fpga_ARADDR_bus[3];
assign \h2f_ARADDR[4]  = hps2fpga_ARADDR_bus[4];
assign \h2f_ARADDR[5]  = hps2fpga_ARADDR_bus[5];
assign \h2f_ARADDR[6]  = hps2fpga_ARADDR_bus[6];
assign \h2f_ARADDR[7]  = hps2fpga_ARADDR_bus[7];
assign \h2f_ARADDR[8]  = hps2fpga_ARADDR_bus[8];
assign \h2f_ARADDR[9]  = hps2fpga_ARADDR_bus[9];
assign \h2f_ARADDR[10]  = hps2fpga_ARADDR_bus[10];
assign \h2f_ARADDR[11]  = hps2fpga_ARADDR_bus[11];
assign \h2f_ARADDR[12]  = hps2fpga_ARADDR_bus[12];
assign \h2f_ARADDR[13]  = hps2fpga_ARADDR_bus[13];
assign \h2f_ARADDR[14]  = hps2fpga_ARADDR_bus[14];
assign \h2f_ARADDR[15]  = hps2fpga_ARADDR_bus[15];
assign \h2f_ARADDR[16]  = hps2fpga_ARADDR_bus[16];
assign \h2f_ARADDR[17]  = hps2fpga_ARADDR_bus[17];
assign \h2f_ARADDR[18]  = hps2fpga_ARADDR_bus[18];
assign \h2f_ARADDR[19]  = hps2fpga_ARADDR_bus[19];
assign \h2f_ARADDR[20]  = hps2fpga_ARADDR_bus[20];
assign \h2f_ARADDR[21]  = hps2fpga_ARADDR_bus[21];
assign \h2f_ARADDR[22]  = hps2fpga_ARADDR_bus[22];
assign \h2f_ARADDR[23]  = hps2fpga_ARADDR_bus[23];
assign \h2f_ARADDR[24]  = hps2fpga_ARADDR_bus[24];
assign \h2f_ARADDR[25]  = hps2fpga_ARADDR_bus[25];
assign \h2f_ARADDR[26]  = hps2fpga_ARADDR_bus[26];
assign \h2f_ARADDR[27]  = hps2fpga_ARADDR_bus[27];
assign \h2f_ARADDR[28]  = hps2fpga_ARADDR_bus[28];
assign \h2f_ARADDR[29]  = hps2fpga_ARADDR_bus[29];

assign \f2sdram~O_BONDING_OUT_10  = f2sdram_BONDING_OUT_1_bus[0];
assign \f2sdram~O_BONDING_OUT_11  = f2sdram_BONDING_OUT_1_bus[1];
assign \f2sdram~O_BONDING_OUT_12  = f2sdram_BONDING_OUT_1_bus[2];
assign \f2sdram~O_BONDING_OUT_13  = f2sdram_BONDING_OUT_1_bus[3];

assign f2h_RDATA[0] = fpga2hps_RDATA_bus[0];
assign f2h_RDATA[1] = fpga2hps_RDATA_bus[1];
assign f2h_RDATA[2] = fpga2hps_RDATA_bus[2];
assign f2h_RDATA[3] = fpga2hps_RDATA_bus[3];
assign f2h_RDATA[4] = fpga2hps_RDATA_bus[4];
assign f2h_RDATA[5] = fpga2hps_RDATA_bus[5];
assign f2h_RDATA[6] = fpga2hps_RDATA_bus[6];
assign f2h_RDATA[7] = fpga2hps_RDATA_bus[7];
assign f2h_RDATA[8] = fpga2hps_RDATA_bus[8];
assign f2h_RDATA[9] = fpga2hps_RDATA_bus[9];
assign f2h_RDATA[10] = fpga2hps_RDATA_bus[10];
assign f2h_RDATA[11] = fpga2hps_RDATA_bus[11];
assign f2h_RDATA[12] = fpga2hps_RDATA_bus[12];
assign f2h_RDATA[13] = fpga2hps_RDATA_bus[13];
assign f2h_RDATA[14] = fpga2hps_RDATA_bus[14];
assign f2h_RDATA[15] = fpga2hps_RDATA_bus[15];
assign f2h_RDATA[16] = fpga2hps_RDATA_bus[16];
assign f2h_RDATA[17] = fpga2hps_RDATA_bus[17];
assign f2h_RDATA[18] = fpga2hps_RDATA_bus[18];
assign f2h_RDATA[19] = fpga2hps_RDATA_bus[19];
assign f2h_RDATA[20] = fpga2hps_RDATA_bus[20];
assign f2h_RDATA[21] = fpga2hps_RDATA_bus[21];
assign f2h_RDATA[22] = fpga2hps_RDATA_bus[22];
assign f2h_RDATA[23] = fpga2hps_RDATA_bus[23];
assign f2h_RDATA[24] = fpga2hps_RDATA_bus[24];
assign f2h_RDATA[25] = fpga2hps_RDATA_bus[25];
assign f2h_RDATA[26] = fpga2hps_RDATA_bus[26];
assign f2h_RDATA[27] = fpga2hps_RDATA_bus[27];
assign f2h_RDATA[28] = fpga2hps_RDATA_bus[28];
assign f2h_RDATA[29] = fpga2hps_RDATA_bus[29];
assign f2h_RDATA[30] = fpga2hps_RDATA_bus[30];
assign f2h_RDATA[31] = fpga2hps_RDATA_bus[31];
assign f2h_RDATA[32] = fpga2hps_RDATA_bus[32];
assign f2h_RDATA[33] = fpga2hps_RDATA_bus[33];
assign f2h_RDATA[34] = fpga2hps_RDATA_bus[34];
assign f2h_RDATA[35] = fpga2hps_RDATA_bus[35];
assign f2h_RDATA[36] = fpga2hps_RDATA_bus[36];
assign f2h_RDATA[37] = fpga2hps_RDATA_bus[37];
assign f2h_RDATA[38] = fpga2hps_RDATA_bus[38];
assign f2h_RDATA[39] = fpga2hps_RDATA_bus[39];
assign f2h_RDATA[40] = fpga2hps_RDATA_bus[40];
assign f2h_RDATA[41] = fpga2hps_RDATA_bus[41];
assign f2h_RDATA[42] = fpga2hps_RDATA_bus[42];
assign f2h_RDATA[43] = fpga2hps_RDATA_bus[43];
assign f2h_RDATA[44] = fpga2hps_RDATA_bus[44];
assign f2h_RDATA[45] = fpga2hps_RDATA_bus[45];
assign f2h_RDATA[46] = fpga2hps_RDATA_bus[46];
assign f2h_RDATA[47] = fpga2hps_RDATA_bus[47];
assign f2h_RDATA[48] = fpga2hps_RDATA_bus[48];
assign f2h_RDATA[49] = fpga2hps_RDATA_bus[49];
assign f2h_RDATA[50] = fpga2hps_RDATA_bus[50];
assign f2h_RDATA[51] = fpga2hps_RDATA_bus[51];
assign f2h_RDATA[52] = fpga2hps_RDATA_bus[52];
assign f2h_RDATA[53] = fpga2hps_RDATA_bus[53];
assign f2h_RDATA[54] = fpga2hps_RDATA_bus[54];
assign f2h_RDATA[55] = fpga2hps_RDATA_bus[55];
assign f2h_RDATA[56] = fpga2hps_RDATA_bus[56];
assign f2h_RDATA[57] = fpga2hps_RDATA_bus[57];
assign f2h_RDATA[58] = fpga2hps_RDATA_bus[58];
assign f2h_RDATA[59] = fpga2hps_RDATA_bus[59];
assign f2h_RDATA[60] = fpga2hps_RDATA_bus[60];
assign f2h_RDATA[61] = fpga2hps_RDATA_bus[61];
assign f2h_RDATA[62] = fpga2hps_RDATA_bus[62];
assign f2h_RDATA[63] = fpga2hps_RDATA_bus[63];

assign h2f_lw_ARADDR[0] = hps2fpga_light_weight_ARADDR_bus[0];
assign h2f_lw_ARADDR[1] = hps2fpga_light_weight_ARADDR_bus[1];
assign h2f_lw_ARADDR[2] = hps2fpga_light_weight_ARADDR_bus[2];
assign h2f_lw_ARADDR[3] = hps2fpga_light_weight_ARADDR_bus[3];
assign h2f_lw_ARADDR[4] = hps2fpga_light_weight_ARADDR_bus[4];
assign h2f_lw_ARADDR[5] = hps2fpga_light_weight_ARADDR_bus[5];
assign \h2f_lw_ARADDR[6]  = hps2fpga_light_weight_ARADDR_bus[6];
assign \h2f_lw_ARADDR[7]  = hps2fpga_light_weight_ARADDR_bus[7];
assign \h2f_lw_ARADDR[8]  = hps2fpga_light_weight_ARADDR_bus[8];
assign \h2f_lw_ARADDR[9]  = hps2fpga_light_weight_ARADDR_bus[9];
assign \h2f_lw_ARADDR[10]  = hps2fpga_light_weight_ARADDR_bus[10];
assign \h2f_lw_ARADDR[11]  = hps2fpga_light_weight_ARADDR_bus[11];
assign \h2f_lw_ARADDR[12]  = hps2fpga_light_weight_ARADDR_bus[12];
assign \h2f_lw_ARADDR[13]  = hps2fpga_light_weight_ARADDR_bus[13];
assign \h2f_lw_ARADDR[14]  = hps2fpga_light_weight_ARADDR_bus[14];
assign \h2f_lw_ARADDR[15]  = hps2fpga_light_weight_ARADDR_bus[15];
assign \h2f_lw_ARADDR[16]  = hps2fpga_light_weight_ARADDR_bus[16];
assign \h2f_lw_ARADDR[17]  = hps2fpga_light_weight_ARADDR_bus[17];
assign \h2f_lw_ARADDR[18]  = hps2fpga_light_weight_ARADDR_bus[18];
assign \h2f_lw_ARADDR[19]  = hps2fpga_light_weight_ARADDR_bus[19];
assign \h2f_lw_ARADDR[20]  = hps2fpga_light_weight_ARADDR_bus[20];

assign h2f_lw_ARBURST[0] = hps2fpga_light_weight_ARBURST_bus[0];
assign h2f_lw_ARBURST[1] = hps2fpga_light_weight_ARBURST_bus[1];

assign h2f_lw_ARID[0] = hps2fpga_light_weight_ARID_bus[0];
assign h2f_lw_ARID[1] = hps2fpga_light_weight_ARID_bus[1];
assign h2f_lw_ARID[2] = hps2fpga_light_weight_ARID_bus[2];
assign h2f_lw_ARID[3] = hps2fpga_light_weight_ARID_bus[3];
assign h2f_lw_ARID[4] = hps2fpga_light_weight_ARID_bus[4];
assign h2f_lw_ARID[5] = hps2fpga_light_weight_ARID_bus[5];
assign h2f_lw_ARID[6] = hps2fpga_light_weight_ARID_bus[6];
assign h2f_lw_ARID[7] = hps2fpga_light_weight_ARID_bus[7];
assign h2f_lw_ARID[8] = hps2fpga_light_weight_ARID_bus[8];
assign h2f_lw_ARID[9] = hps2fpga_light_weight_ARID_bus[9];
assign h2f_lw_ARID[10] = hps2fpga_light_weight_ARID_bus[10];
assign h2f_lw_ARID[11] = hps2fpga_light_weight_ARID_bus[11];

assign h2f_lw_ARLEN[0] = hps2fpga_light_weight_ARLEN_bus[0];
assign h2f_lw_ARLEN[1] = hps2fpga_light_weight_ARLEN_bus[1];
assign h2f_lw_ARLEN[2] = hps2fpga_light_weight_ARLEN_bus[2];
assign h2f_lw_ARLEN[3] = hps2fpga_light_weight_ARLEN_bus[3];

assign h2f_lw_ARSIZE[0] = hps2fpga_light_weight_ARSIZE_bus[0];
assign h2f_lw_ARSIZE[1] = hps2fpga_light_weight_ARSIZE_bus[1];
assign h2f_lw_ARSIZE[2] = hps2fpga_light_weight_ARSIZE_bus[2];

assign h2f_lw_AWADDR[0] = hps2fpga_light_weight_AWADDR_bus[0];
assign h2f_lw_AWADDR[1] = hps2fpga_light_weight_AWADDR_bus[1];
assign h2f_lw_AWADDR[2] = hps2fpga_light_weight_AWADDR_bus[2];
assign h2f_lw_AWADDR[3] = hps2fpga_light_weight_AWADDR_bus[3];
assign h2f_lw_AWADDR[4] = hps2fpga_light_weight_AWADDR_bus[4];
assign h2f_lw_AWADDR[5] = hps2fpga_light_weight_AWADDR_bus[5];

assign h2f_lw_AWBURST[0] = hps2fpga_light_weight_AWBURST_bus[0];
assign h2f_lw_AWBURST[1] = hps2fpga_light_weight_AWBURST_bus[1];

assign h2f_lw_AWID[0] = hps2fpga_light_weight_AWID_bus[0];
assign h2f_lw_AWID[1] = hps2fpga_light_weight_AWID_bus[1];
assign h2f_lw_AWID[2] = hps2fpga_light_weight_AWID_bus[2];
assign h2f_lw_AWID[3] = hps2fpga_light_weight_AWID_bus[3];
assign h2f_lw_AWID[4] = hps2fpga_light_weight_AWID_bus[4];
assign h2f_lw_AWID[5] = hps2fpga_light_weight_AWID_bus[5];
assign h2f_lw_AWID[6] = hps2fpga_light_weight_AWID_bus[6];
assign h2f_lw_AWID[7] = hps2fpga_light_weight_AWID_bus[7];
assign h2f_lw_AWID[8] = hps2fpga_light_weight_AWID_bus[8];
assign h2f_lw_AWID[9] = hps2fpga_light_weight_AWID_bus[9];
assign h2f_lw_AWID[10] = hps2fpga_light_weight_AWID_bus[10];
assign h2f_lw_AWID[11] = hps2fpga_light_weight_AWID_bus[11];

assign h2f_lw_AWLEN[0] = hps2fpga_light_weight_AWLEN_bus[0];
assign h2f_lw_AWLEN[1] = hps2fpga_light_weight_AWLEN_bus[1];
assign h2f_lw_AWLEN[2] = hps2fpga_light_weight_AWLEN_bus[2];
assign h2f_lw_AWLEN[3] = hps2fpga_light_weight_AWLEN_bus[3];

assign h2f_lw_AWSIZE[0] = hps2fpga_light_weight_AWSIZE_bus[0];
assign h2f_lw_AWSIZE[1] = hps2fpga_light_weight_AWSIZE_bus[1];
assign h2f_lw_AWSIZE[2] = hps2fpga_light_weight_AWSIZE_bus[2];

assign h2f_lw_WDATA[0] = hps2fpga_light_weight_WDATA_bus[0];
assign h2f_lw_WDATA[1] = hps2fpga_light_weight_WDATA_bus[1];
assign h2f_lw_WDATA[2] = hps2fpga_light_weight_WDATA_bus[2];
assign h2f_lw_WDATA[3] = hps2fpga_light_weight_WDATA_bus[3];
assign h2f_lw_WDATA[4] = hps2fpga_light_weight_WDATA_bus[4];
assign h2f_lw_WDATA[5] = hps2fpga_light_weight_WDATA_bus[5];
assign h2f_lw_WDATA[6] = hps2fpga_light_weight_WDATA_bus[6];
assign h2f_lw_WDATA[7] = hps2fpga_light_weight_WDATA_bus[7];
assign h2f_lw_WDATA[8] = hps2fpga_light_weight_WDATA_bus[8];
assign h2f_lw_WDATA[9] = hps2fpga_light_weight_WDATA_bus[9];
assign h2f_lw_WDATA[10] = hps2fpga_light_weight_WDATA_bus[10];
assign h2f_lw_WDATA[11] = hps2fpga_light_weight_WDATA_bus[11];
assign h2f_lw_WDATA[12] = hps2fpga_light_weight_WDATA_bus[12];
assign h2f_lw_WDATA[13] = hps2fpga_light_weight_WDATA_bus[13];
assign h2f_lw_WDATA[14] = hps2fpga_light_weight_WDATA_bus[14];
assign h2f_lw_WDATA[15] = hps2fpga_light_weight_WDATA_bus[15];
assign h2f_lw_WDATA[16] = hps2fpga_light_weight_WDATA_bus[16];
assign h2f_lw_WDATA[17] = hps2fpga_light_weight_WDATA_bus[17];
assign h2f_lw_WDATA[18] = hps2fpga_light_weight_WDATA_bus[18];
assign h2f_lw_WDATA[19] = hps2fpga_light_weight_WDATA_bus[19];
assign h2f_lw_WDATA[20] = hps2fpga_light_weight_WDATA_bus[20];
assign h2f_lw_WDATA[21] = hps2fpga_light_weight_WDATA_bus[21];
assign h2f_lw_WDATA[22] = hps2fpga_light_weight_WDATA_bus[22];
assign h2f_lw_WDATA[23] = hps2fpga_light_weight_WDATA_bus[23];
assign h2f_lw_WDATA[24] = hps2fpga_light_weight_WDATA_bus[24];
assign h2f_lw_WDATA[25] = hps2fpga_light_weight_WDATA_bus[25];
assign h2f_lw_WDATA[26] = hps2fpga_light_weight_WDATA_bus[26];
assign h2f_lw_WDATA[27] = hps2fpga_light_weight_WDATA_bus[27];
assign h2f_lw_WDATA[28] = hps2fpga_light_weight_WDATA_bus[28];
assign h2f_lw_WDATA[29] = hps2fpga_light_weight_WDATA_bus[29];
assign h2f_lw_WDATA[30] = hps2fpga_light_weight_WDATA_bus[30];
assign h2f_lw_WDATA[31] = hps2fpga_light_weight_WDATA_bus[31];

assign h2f_lw_WSTRB[0] = hps2fpga_light_weight_WSTRB_bus[0];
assign h2f_lw_WSTRB[1] = hps2fpga_light_weight_WSTRB_bus[1];
assign h2f_lw_WSTRB[2] = hps2fpga_light_weight_WSTRB_bus[2];
assign h2f_lw_WSTRB[3] = hps2fpga_light_weight_WSTRB_bus[3];

cyclonev_hps_interface_clocks_resets clocks_resets(
	.f2h_cold_rst_req_n(vcc),
	.f2h_dbg_rst_req_n(vcc),
	.f2h_pending_rst_ack(vcc),
	.f2h_periph_ref_clk(gnd),
	.f2h_sdram_ref_clk(gnd),
	.f2h_warm_rst_req_n(vcc),
	.ptp_ref_clk(gnd),
	.h2f_cold_rst_n(\clocks_resets~h2f_cold_rst_n ),
	.h2f_pending_rst_req_n(),
	.h2f_rst_n(h2f_rst_n[0]),
	.h2f_user0_clk(),
	.h2f_user1_clk(),
	.h2f_user2_clk());
defparam clocks_resets.h2f_user0_clk_freq = 100;
defparam clocks_resets.h2f_user1_clk_freq = 100;
defparam clocks_resets.h2f_user2_clk_freq = 100;

cyclonev_hps_interface_fpga2hps fpga2hps(
	.arvalid(f2h_ARVALID[0]),
	.awvalid(f2h_AWVALID[0]),
	.bready(f2h_BREADY[0]),
	.clk(h2f_lw_axi_clk[0]),
	.rready(f2h_RVALID[0]),
	.wlast(f2h_AWSIZE[1]),
	.wvalid(f2h_WVALID[0]),
	.araddr({f2h_ARADDR[31],f2h_ARADDR[30],f2h_ARADDR[29],f2h_ARADDR[28],f2h_ARADDR[27],f2h_ARADDR[26],f2h_ARADDR[25],f2h_ARADDR[24],f2h_ARADDR[23],f2h_ARADDR[22],f2h_ARADDR[21],f2h_ARADDR[20],f2h_ARADDR[19],f2h_ARADDR[18],f2h_ARADDR[17],f2h_ARADDR[16],f2h_ARADDR[15],f2h_ARADDR[14],f2h_ARADDR[13],f2h_ARADDR[12],f2h_ARADDR[11],f2h_ARADDR[10],f2h_ARADDR[9],f2h_ARADDR[8],f2h_ARADDR[7],
f2h_ARADDR[6],f2h_ARADDR[5],f2h_ARADDR[4],f2h_ARADDR[3],f2h_ARADDR[2],gnd,gnd}),
	.arburst({gnd,f2h_ARSIZE[1]}),
	.arcache({gnd,gnd,gnd,gnd}),
	.arid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arlen({gnd,gnd,gnd,gnd}),
	.arlock({gnd,gnd}),
	.arprot({gnd,f2h_ARSIZE[1],gnd}),
	.arsize({gnd,f2h_ARSIZE[1],gnd}),
	.aruser({gnd,gnd,gnd,gnd,gnd}),
	.awaddr({f2h_AWADDR[31],f2h_AWADDR[30],f2h_AWADDR[29],f2h_AWADDR[28],f2h_AWADDR[27],f2h_AWADDR[26],f2h_AWADDR[25],f2h_AWADDR[24],f2h_AWADDR[23],f2h_AWADDR[22],f2h_AWADDR[21],f2h_AWADDR[20],f2h_AWADDR[19],f2h_AWADDR[18],f2h_AWADDR[17],f2h_AWADDR[16],f2h_AWADDR[15],f2h_AWADDR[14],f2h_AWADDR[13],f2h_AWADDR[12],f2h_AWADDR[11],f2h_AWADDR[10],f2h_AWADDR[9],f2h_AWADDR[8],f2h_AWADDR[7],
f2h_AWADDR[6],f2h_AWADDR[5],f2h_AWADDR[4],f2h_AWADDR[3],f2h_AWADDR[2],gnd,gnd}),
	.awburst({gnd,f2h_AWSIZE[1]}),
	.awcache({gnd,gnd,gnd,gnd}),
	.awid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awlen({!f2h_AWSIZE[1],!f2h_AWSIZE[1],!f2h_AWSIZE[1],!f2h_AWSIZE[1]}),
	.awlock({gnd,gnd}),
	.awprot({gnd,f2h_AWSIZE[1],gnd}),
	.awsize({gnd,f2h_AWSIZE[1],gnd}),
	.awuser({gnd,gnd,gnd,gnd,gnd}),
	.port_size_config({gnd,vcc}),
	.wdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_WDATA[63],f2h_WDATA[62],f2h_WDATA[61],f2h_WDATA[60],f2h_WDATA[59],f2h_WDATA[58],f2h_WDATA[57],
f2h_WDATA[56],f2h_WDATA[55],f2h_WDATA[54],f2h_WDATA[53],f2h_WDATA[52],f2h_WDATA[51],f2h_WDATA[50],f2h_WDATA[49],f2h_WDATA[48],f2h_WDATA[47],f2h_WDATA[46],f2h_WDATA[45],f2h_WDATA[44],f2h_WDATA[43],f2h_WDATA[42],f2h_WDATA[41],f2h_WDATA[40],f2h_WDATA[39],f2h_WDATA[38],f2h_WDATA[37],f2h_WDATA[36],f2h_WDATA[35],f2h_WDATA[34],f2h_WDATA[33],f2h_WDATA[32],f2h_WDATA[31],f2h_WDATA[30],f2h_WDATA[29],
f2h_WDATA[28],f2h_WDATA[27],f2h_WDATA[26],f2h_WDATA[25],f2h_WDATA[24],f2h_WDATA[23],f2h_WDATA[22],f2h_WDATA[21],f2h_WDATA[20],f2h_WDATA[19],f2h_WDATA[18],f2h_WDATA[17],f2h_WDATA[16],f2h_WDATA[15],f2h_WDATA[14],f2h_WDATA[13],f2h_WDATA[12],f2h_WDATA[11],f2h_WDATA[10],f2h_WDATA[9],f2h_WDATA[8],f2h_WDATA[7],f2h_WDATA[6],f2h_WDATA[5],f2h_WDATA[4],f2h_WDATA[3],f2h_WDATA[2],f2h_WDATA[1],
f2h_WDATA[0]}),
	.wid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wstrb({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_WSTRB[7],f2h_WSTRB[6],f2h_WSTRB[5],f2h_WSTRB[4],f2h_WSTRB[3],f2h_WSTRB[2],f2h_WSTRB[1],f2h_WSTRB[0]}),
	.arready(f2h_ARREADY[0]),
	.awready(f2h_AWREADY[0]),
	.bvalid(f2h_BVALID[0]),
	.rlast(),
	.rvalid(f2h_RVALID[0]),
	.wready(f2h_WREADY[0]),
	.bid(),
	.bresp(),
	.rdata(fpga2hps_RDATA_bus),
	.rid(),
	.rresp());
defparam fpga2hps.data_width = 32;

cyclonev_hps_interface_hps2fpga_light_weight hps2fpga_light_weight(
	.arready(h2f_lw_ARREADY[0]),
	.awready(h2f_lw_AWREADY[0]),
	.bvalid(h2f_lw_BVALID[0]),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(h2f_lw_RLAST[0]),
	.rvalid(h2f_lw_RVALID[0]),
	.wready(h2f_lw_WREADY[0]),
	.bid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.bresp({gnd,gnd}),
	.rdata({h2f_lw_RDATA[31],h2f_lw_RDATA[30],h2f_lw_RDATA[29],h2f_lw_RDATA[28],h2f_lw_RDATA[27],h2f_lw_RDATA[26],h2f_lw_RDATA[25],h2f_lw_RDATA[24],h2f_lw_RDATA[23],h2f_lw_RDATA[22],h2f_lw_RDATA[21],h2f_lw_RDATA[20],h2f_lw_RDATA[19],h2f_lw_RDATA[18],h2f_lw_RDATA[17],h2f_lw_RDATA[16],h2f_lw_RDATA[15],h2f_lw_RDATA[14],h2f_lw_RDATA[13],h2f_lw_RDATA[12],h2f_lw_RDATA[11],
h2f_lw_RDATA[10],h2f_lw_RDATA[9],h2f_lw_RDATA[8],h2f_lw_RDATA[7],h2f_lw_RDATA[6],h2f_lw_RDATA[5],h2f_lw_RDATA[4],h2f_lw_RDATA[3],h2f_lw_RDATA[2],h2f_lw_RDATA[1],h2f_lw_RDATA[0]}),
	.rid({h2f_lw_RID[11],h2f_lw_RID[10],h2f_lw_RID[9],h2f_lw_RID[8],h2f_lw_RID[7],h2f_lw_RID[6],h2f_lw_RID[5],h2f_lw_RID[4],h2f_lw_RID[3],h2f_lw_RID[2],h2f_lw_RID[1],h2f_lw_RID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_lw_ARVALID[0]),
	.awvalid(h2f_lw_AWVALID[0]),
	.bready(h2f_lw_BREADY[0]),
	.rready(h2f_lw_RREADY[0]),
	.wlast(h2f_lw_WLAST[0]),
	.wvalid(h2f_lw_WVALID[0]),
	.araddr(hps2fpga_light_weight_ARADDR_bus),
	.arburst(hps2fpga_light_weight_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_light_weight_ARID_bus),
	.arlen(hps2fpga_light_weight_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_light_weight_ARSIZE_bus),
	.awaddr(hps2fpga_light_weight_AWADDR_bus),
	.awburst(hps2fpga_light_weight_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_light_weight_AWID_bus),
	.awlen(hps2fpga_light_weight_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_light_weight_AWSIZE_bus),
	.wdata(hps2fpga_light_weight_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_light_weight_WSTRB_bus));

cyclonev_hps_interface_dbg_apb debug_apb(
	.p_slv_err(gnd),
	.p_ready(gnd),
	.p_clk(gnd),
	.p_clk_en(gnd),
	.dbg_apb_disable(gnd),
	.p_rdata(32'b00000000000000000000000000000000),
	.p_addr_31(\debug_apb~O_P_ADDR_31 ),
	.p_write(),
	.p_sel(),
	.p_enable(),
	.p_reset_n(),
	.p_addr(),
	.p_wdata());
defparam debug_apb.dummy_param = 256;

cyclonev_hps_interface_tpiu_trace tpiu(
	.traceclk_ctl(vcc),
	.traceclkin(gnd),
	.traceclk(),
	.trace_data(tpiu_TRACE_DATA_bus));

cyclonev_hps_interface_boot_from_fpga boot_from_fpga(
	.boot_from_fpga_on_failure(gnd),
	.boot_from_fpga_ready(gnd),
	.bsel_en(gnd),
	.csel_en(gnd),
	.bsel({gnd,gnd,vcc}),
	.csel({gnd,vcc}),
	.fake_dout(\boot_from_fpga~fake_dout ));

cyclonev_hps_interface_hps2fpga hps2fpga(
	.arready(gnd),
	.awready(gnd),
	.bvalid(gnd),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(gnd),
	.rvalid(gnd),
	.wready(gnd),
	.bid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.bresp({gnd,gnd}),
	.port_size_config({vcc,gnd}),
	.rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rresp({gnd,gnd}),
	.arvalid(),
	.awvalid(),
	.bready(),
	.rready(),
	.wlast(),
	.wvalid(),
	.araddr(hps2fpga_ARADDR_bus),
	.arburst(),
	.arcache(),
	.arid(),
	.arlen(),
	.arlock(),
	.arprot(),
	.arsize(),
	.awaddr(),
	.awburst(),
	.awcache(),
	.awid(),
	.awlen(),
	.awlock(),
	.awprot(),
	.awsize(),
	.wdata(),
	.wid(),
	.wstrb());
defparam hps2fpga.data_width = 32;

cyclonev_hps_interface_fpga2sdram f2sdram(
	.cmd_port_clk_0(gnd),
	.cmd_port_clk_1(gnd),
	.cmd_port_clk_2(gnd),
	.cmd_port_clk_3(gnd),
	.cmd_port_clk_4(gnd),
	.cmd_port_clk_5(gnd),
	.cmd_valid_0(gnd),
	.cmd_valid_1(gnd),
	.cmd_valid_2(gnd),
	.cmd_valid_3(gnd),
	.cmd_valid_4(gnd),
	.cmd_valid_5(gnd),
	.rd_clk_0(gnd),
	.rd_clk_1(gnd),
	.rd_clk_2(gnd),
	.rd_clk_3(gnd),
	.rd_ready_0(gnd),
	.rd_ready_1(gnd),
	.rd_ready_2(gnd),
	.rd_ready_3(gnd),
	.wr_clk_0(gnd),
	.wr_clk_1(gnd),
	.wr_clk_2(gnd),
	.wr_clk_3(gnd),
	.wr_valid_0(gnd),
	.wr_valid_1(gnd),
	.wr_valid_2(gnd),
	.wr_valid_3(gnd),
	.wrack_ready_0(gnd),
	.wrack_ready_1(gnd),
	.wrack_ready_2(gnd),
	.wrack_ready_3(gnd),
	.wrack_ready_4(gnd),
	.wrack_ready_5(gnd),
	.cfg_axi_mm_select({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_rfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_type({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_wfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_port_width({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_rfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_wfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_data_0(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_1(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_2(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_3(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_4(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_5(60'b000000000000000000000000000000000000000000000000000000000000),
	.wr_data_0(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_1(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_2(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_3(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.cmd_ready_0(),
	.cmd_ready_1(),
	.cmd_ready_2(),
	.cmd_ready_3(),
	.cmd_ready_4(),
	.cmd_ready_5(),
	.rd_valid_0(),
	.rd_valid_1(),
	.rd_valid_2(),
	.rd_valid_3(),
	.wr_ready_0(),
	.wr_ready_1(),
	.wr_ready_2(),
	.wr_ready_3(),
	.wrack_valid_0(),
	.wrack_valid_1(),
	.wrack_valid_2(),
	.wrack_valid_3(),
	.wrack_valid_4(),
	.wrack_valid_5(),
	.bonding_out_1(f2sdram_BONDING_OUT_1_bus),
	.bonding_out_2(),
	.rd_data_0(),
	.rd_data_1(),
	.rd_data_2(),
	.rd_data_3(),
	.wrack_data_0(),
	.wrack_data_1(),
	.wrack_data_2(),
	.wrack_data_3(),
	.wrack_data_4(),
	.wrack_data_5());

cyclonev_hps_interface_interrupts interrupts(
	.irq({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_irq_p0[31],f2h_irq_p0[30],f2h_irq_p0[29],f2h_irq_p0[28],f2h_irq_p0[27],f2h_irq_p0[26],f2h_irq_p0[25],f2h_irq_p0[24],f2h_irq_p0[23],f2h_irq_p0[22],f2h_irq_p0[21],f2h_irq_p0[20],f2h_irq_p0[19],f2h_irq_p0[18],f2h_irq_p0[17],f2h_irq_p0[16],
f2h_irq_p0[15],f2h_irq_p0[14],f2h_irq_p0[13],f2h_irq_p0[12],f2h_irq_p0[11],f2h_irq_p0[10],f2h_irq_p0[9],f2h_irq_p0[8],f2h_irq_p0[7],f2h_irq_p0[6],f2h_irq_p0[5],f2h_irq_p0[4],f2h_irq_p0[3],f2h_irq_p0[2],f2h_irq_p0[1],f2h_irq_p0[0]}),
	.fake_dout(\interrupts~fake_dout ),
	.h2f_can0_irq(),
	.h2f_can1_irq(),
	.h2f_clkmgr_irq(),
	.h2f_cti_irq0_n(),
	.h2f_cti_irq1_n(),
	.h2f_dma_abort_irq(),
	.h2f_dma_irq0(),
	.h2f_dma_irq1(),
	.h2f_dma_irq2(),
	.h2f_dma_irq3(),
	.h2f_dma_irq4(),
	.h2f_dma_irq5(),
	.h2f_dma_irq6(),
	.h2f_dma_irq7(),
	.h2f_emac0_irq(),
	.h2f_emac1_irq(),
	.h2f_fpga_man_irq(),
	.h2f_gpio0_irq(),
	.h2f_gpio1_irq(),
	.h2f_gpio2_irq(),
	.h2f_i2c0_irq(),
	.h2f_i2c1_irq(),
	.h2f_i2c_emac0_irq(),
	.h2f_i2c_emac1_irq(),
	.h2f_l4sp0_irq(),
	.h2f_l4sp1_irq(),
	.h2f_mpuwakeup_irq(),
	.h2f_nand_irq(),
	.h2f_osc0_irq(),
	.h2f_osc1_irq(),
	.h2f_qspi_irq(),
	.h2f_sdmmc_irq(),
	.h2f_spi0_irq(),
	.h2f_spi1_irq(),
	.h2f_spi2_irq(),
	.h2f_spi3_irq(),
	.h2f_uart0_irq(),
	.h2f_uart1_irq(),
	.h2f_usb0_irq(),
	.h2f_usb1_irq(),
	.h2f_wdog0_irq(),
	.h2f_wdog1_irq());

endmodule

module Computer_System_Computer_System_ARM_A9_HPS_hps_io (
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim1_inst,
	spim1_inst1,
	intermediate_36,
	intermediate_37,
	uart0_inst,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	intermediate_42,
	intermediate_43,
	intermediate_44,
	intermediate_46,
	intermediate_48,
	intermediate_50,
	intermediate_52,
	intermediate_54,
	intermediate_45,
	intermediate_47,
	intermediate_49,
	intermediate_51,
	intermediate_53,
	intermediate_55,
	intermediate_56,
	intermediate_57,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO35_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO41_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO53_0,
	hps_io_gpio_inst_GPIO54_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	uart0_inst;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	intermediate_42;
output 	intermediate_43;
output 	intermediate_44;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_50;
output 	intermediate_52;
output 	intermediate_54;
output 	intermediate_45;
output 	intermediate_47;
output 	intermediate_49;
output 	intermediate_51;
output 	intermediate_53;
output 	intermediate_55;
output 	intermediate_56;
output 	intermediate_57;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO35_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO41_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO53_0;
input 	hps_io_gpio_inst_GPIO54_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_ARM_A9_HPS_hps_io_border border(
	.hps_io_emac1_inst_TX_CLK({emac1_inst}),
	.hps_io_emac1_inst_TX_CTL({emac1_inst1}),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.hps_io_emac1_inst_MDC({emac1_inst2}),
	.hps_io_emac1_inst_TXD0({emac1_inst3}),
	.hps_io_emac1_inst_TXD1({emac1_inst4}),
	.hps_io_emac1_inst_TXD2({emac1_inst5}),
	.hps_io_emac1_inst_TXD3({emac1_inst6}),
	.hps_io_qspi_inst_CLK({qspi_inst}),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.hps_io_qspi_inst_SS0({qspi_inst1}),
	.hps_io_sdio_inst_CLK({sdio_inst}),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.hps_io_usb1_inst_STP({usb1_inst}),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.hps_io_spim1_inst_CLK({spim1_inst}),
	.hps_io_spim1_inst_SS0({spim1_inst1}),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.hps_io_uart0_inst_TX({uart0_inst}),
	.intermediate_39(intermediate_39),
	.intermediate_38(intermediate_38),
	.intermediate_41(intermediate_41),
	.intermediate_40(intermediate_40),
	.intermediate_42(intermediate_42),
	.intermediate_43(intermediate_43),
	.intermediate_44(intermediate_44),
	.intermediate_46(intermediate_46),
	.intermediate_48(intermediate_48),
	.intermediate_50(intermediate_50),
	.intermediate_52(intermediate_52),
	.intermediate_54(intermediate_54),
	.intermediate_45(intermediate_45),
	.intermediate_47(intermediate_47),
	.intermediate_49(intermediate_49),
	.intermediate_51(intermediate_51),
	.intermediate_53(intermediate_53),
	.intermediate_55(intermediate_55),
	.intermediate_56(intermediate_56),
	.intermediate_57(intermediate_57),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_i2c0_inst_SDA_0(hps_io_i2c0_inst_SDA_0),
	.hps_io_i2c0_inst_SCL_0(hps_io_i2c0_inst_SCL_0),
	.hps_io_i2c1_inst_SDA_0(hps_io_i2c1_inst_SDA_0),
	.hps_io_i2c1_inst_SCL_0(hps_io_i2c1_inst_SCL_0),
	.hps_io_gpio_inst_GPIO09_0(hps_io_gpio_inst_GPIO09_0),
	.hps_io_gpio_inst_GPIO35_0(hps_io_gpio_inst_GPIO35_0),
	.hps_io_gpio_inst_GPIO40_0(hps_io_gpio_inst_GPIO40_0),
	.hps_io_gpio_inst_GPIO41_0(hps_io_gpio_inst_GPIO41_0),
	.hps_io_gpio_inst_GPIO48_0(hps_io_gpio_inst_GPIO48_0),
	.hps_io_gpio_inst_GPIO53_0(hps_io_gpio_inst_GPIO53_0),
	.hps_io_gpio_inst_GPIO54_0(hps_io_gpio_inst_GPIO54_0),
	.hps_io_gpio_inst_GPIO61_0(hps_io_gpio_inst_GPIO61_0),
	.hps_io_emac1_inst_RXD0({hps_io_hps_io_emac1_inst_RXD0}),
	.hps_io_emac1_inst_RXD1({hps_io_hps_io_emac1_inst_RXD1}),
	.hps_io_emac1_inst_RXD2({hps_io_hps_io_emac1_inst_RXD2}),
	.hps_io_emac1_inst_RXD3({hps_io_hps_io_emac1_inst_RXD3}),
	.hps_io_emac1_inst_RX_CLK({hps_io_hps_io_emac1_inst_RX_CLK}),
	.hps_io_emac1_inst_RX_CTL({hps_io_hps_io_emac1_inst_RX_CTL}),
	.hps_io_spim1_inst_MISO({hps_io_hps_io_spim1_inst_MISO}),
	.hps_io_uart0_inst_RX({hps_io_hps_io_uart0_inst_RX}),
	.hps_io_usb1_inst_CLK({hps_io_hps_io_usb1_inst_CLK}),
	.hps_io_usb1_inst_DIR({hps_io_hps_io_usb1_inst_DIR}),
	.hps_io_usb1_inst_NXT({hps_io_hps_io_usb1_inst_NXT}),
	.memory_oct_rzqin(memory_oct_rzqin));

endmodule

module Computer_System_Computer_System_ARM_A9_HPS_hps_io_border (
	hps_io_emac1_inst_TX_CLK,
	hps_io_emac1_inst_TX_CTL,
	intermediate_0,
	intermediate_1,
	hps_io_emac1_inst_MDC,
	hps_io_emac1_inst_TXD0,
	hps_io_emac1_inst_TXD1,
	hps_io_emac1_inst_TXD2,
	hps_io_emac1_inst_TXD3,
	hps_io_qspi_inst_CLK,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	hps_io_qspi_inst_SS0,
	hps_io_sdio_inst_CLK,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	hps_io_usb1_inst_STP,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	hps_io_spim1_inst_CLK,
	hps_io_spim1_inst_SS0,
	intermediate_36,
	intermediate_37,
	hps_io_uart0_inst_TX,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	intermediate_42,
	intermediate_43,
	intermediate_44,
	intermediate_46,
	intermediate_48,
	intermediate_50,
	intermediate_52,
	intermediate_54,
	intermediate_45,
	intermediate_47,
	intermediate_49,
	intermediate_51,
	intermediate_53,
	intermediate_55,
	intermediate_56,
	intermediate_57,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO35_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO41_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO53_0,
	hps_io_gpio_inst_GPIO54_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_emac1_inst_RXD0,
	hps_io_emac1_inst_RXD1,
	hps_io_emac1_inst_RXD2,
	hps_io_emac1_inst_RXD3,
	hps_io_emac1_inst_RX_CLK,
	hps_io_emac1_inst_RX_CTL,
	hps_io_spim1_inst_MISO,
	hps_io_uart0_inst_RX,
	hps_io_usb1_inst_CLK,
	hps_io_usb1_inst_DIR,
	hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[0:0] hps_io_emac1_inst_TX_CLK;
output 	[0:0] hps_io_emac1_inst_TX_CTL;
output 	intermediate_0;
output 	intermediate_1;
output 	[0:0] hps_io_emac1_inst_MDC;
output 	[0:0] hps_io_emac1_inst_TXD0;
output 	[0:0] hps_io_emac1_inst_TXD1;
output 	[0:0] hps_io_emac1_inst_TXD2;
output 	[0:0] hps_io_emac1_inst_TXD3;
output 	[0:0] hps_io_qspi_inst_CLK;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	[0:0] hps_io_qspi_inst_SS0;
output 	[0:0] hps_io_sdio_inst_CLK;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	[0:0] hps_io_usb1_inst_STP;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	[0:0] hps_io_spim1_inst_CLK;
output 	[0:0] hps_io_spim1_inst_SS0;
output 	intermediate_36;
output 	intermediate_37;
output 	[0:0] hps_io_uart0_inst_TX;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	intermediate_42;
output 	intermediate_43;
output 	intermediate_44;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_50;
output 	intermediate_52;
output 	intermediate_54;
output 	intermediate_45;
output 	intermediate_47;
output 	intermediate_49;
output 	intermediate_51;
output 	intermediate_53;
output 	intermediate_55;
output 	intermediate_56;
output 	intermediate_57;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO35_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO41_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO53_0;
input 	hps_io_gpio_inst_GPIO54_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	[0:0] hps_io_emac1_inst_RXD0;
input 	[0:0] hps_io_emac1_inst_RXD1;
input 	[0:0] hps_io_emac1_inst_RXD2;
input 	[0:0] hps_io_emac1_inst_RXD3;
input 	[0:0] hps_io_emac1_inst_RX_CLK;
input 	[0:0] hps_io_emac1_inst_RX_CTL;
input 	[0:0] hps_io_spim1_inst_MISO;
input 	[0:0] hps_io_uart0_inst_RX;
input 	[0:0] hps_io_usb1_inst_CLK;
input 	[0:0] hps_io_usb1_inst_DIR;
input 	[0:0] hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdio_inst~O_SDMMC_PWR_EN ;
wire \uart0_inst~UARTRTSN ;
wire \gpio_inst~LOANIO0_I0 ;
wire \gpio_inst~LOANIO0_I1 ;
wire \gpio_inst~LOANIO0_I2 ;
wire \gpio_inst~LOANIO0_I3 ;
wire \gpio_inst~LOANIO0_I4 ;
wire \gpio_inst~LOANIO0_I5 ;
wire \gpio_inst~LOANIO0_I6 ;
wire \gpio_inst~LOANIO0_I7 ;
wire \gpio_inst~LOANIO0_I8 ;
wire \gpio_inst~LOANIO0_I9 ;
wire \gpio_inst~LOANIO0_I10 ;
wire \gpio_inst~LOANIO0_I11 ;
wire \gpio_inst~LOANIO0_I12 ;
wire \gpio_inst~LOANIO0_I13 ;
wire \gpio_inst~LOANIO0_I14 ;
wire \gpio_inst~LOANIO0_I15 ;
wire \gpio_inst~LOANIO0_I16 ;
wire \gpio_inst~LOANIO0_I17 ;
wire \gpio_inst~LOANIO0_I18 ;
wire \gpio_inst~LOANIO0_I19 ;
wire \gpio_inst~LOANIO0_I20 ;
wire \gpio_inst~LOANIO0_I21 ;
wire \gpio_inst~LOANIO0_I22 ;
wire \gpio_inst~LOANIO0_I23 ;
wire \gpio_inst~LOANIO0_I24 ;
wire \gpio_inst~LOANIO0_I25 ;
wire \gpio_inst~LOANIO0_I26 ;
wire \gpio_inst~LOANIO0_I27 ;
wire \gpio_inst~LOANIO0_I28 ;
wire \~GND~combout ;

wire [3:0] emac1_inst_EMAC_PHY_TXD_bus;
wire [3:0] qspi_inst_QSPI_SS_N_bus;
wire [3:0] qspi_inst_QSPI_MO_EN_N_bus;
wire [7:0] sdio_inst_SDMMC_DATA_OE_bus;
wire [7:0] sdio_inst_SDMMC_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_OE_bus;
wire [28:0] gpio_inst_GPIO1_PORTA_O_bus;
wire [28:0] gpio_inst_GPIO0_PORTA_OE_bus;
wire [12:0] gpio_inst_GPIO2_PORTA_O_bus;
wire [28:0] gpio_inst_GPIO0_PORTA_O_bus;
wire [12:0] gpio_inst_GPIO2_PORTA_OE_bus;
wire [28:0] gpio_inst_GPIO1_PORTA_OE_bus;
wire [28:0] gpio_inst_LOANIO0_I_bus;

assign hps_io_emac1_inst_TXD0[0] = emac1_inst_EMAC_PHY_TXD_bus[0];
assign hps_io_emac1_inst_TXD1[0] = emac1_inst_EMAC_PHY_TXD_bus[1];
assign hps_io_emac1_inst_TXD2[0] = emac1_inst_EMAC_PHY_TXD_bus[2];
assign hps_io_emac1_inst_TXD3[0] = emac1_inst_EMAC_PHY_TXD_bus[3];

assign hps_io_qspi_inst_SS0[0] = qspi_inst_QSPI_SS_N_bus[0];

assign intermediate_3 = qspi_inst_QSPI_MO_EN_N_bus[0];
assign intermediate_5 = qspi_inst_QSPI_MO_EN_N_bus[1];
assign intermediate_7 = qspi_inst_QSPI_MO_EN_N_bus[2];
assign intermediate_9 = qspi_inst_QSPI_MO_EN_N_bus[3];

assign intermediate_13 = sdio_inst_SDMMC_DATA_OE_bus[0];
assign intermediate_15 = sdio_inst_SDMMC_DATA_OE_bus[1];
assign intermediate_17 = sdio_inst_SDMMC_DATA_OE_bus[2];
assign intermediate_19 = sdio_inst_SDMMC_DATA_OE_bus[3];

assign intermediate_12 = sdio_inst_SDMMC_DATA_O_bus[0];
assign intermediate_14 = sdio_inst_SDMMC_DATA_O_bus[1];
assign intermediate_16 = sdio_inst_SDMMC_DATA_O_bus[2];
assign intermediate_18 = sdio_inst_SDMMC_DATA_O_bus[3];

assign intermediate_20 = usb1_inst_USB_ULPI_DATA_O_bus[0];
assign intermediate_22 = usb1_inst_USB_ULPI_DATA_O_bus[1];
assign intermediate_24 = usb1_inst_USB_ULPI_DATA_O_bus[2];
assign intermediate_26 = usb1_inst_USB_ULPI_DATA_O_bus[3];
assign intermediate_28 = usb1_inst_USB_ULPI_DATA_O_bus[4];
assign intermediate_30 = usb1_inst_USB_ULPI_DATA_O_bus[5];
assign intermediate_32 = usb1_inst_USB_ULPI_DATA_O_bus[6];
assign intermediate_34 = usb1_inst_USB_ULPI_DATA_O_bus[7];

assign intermediate_21 = usb1_inst_USB_ULPI_DATA_OE_bus[0];
assign intermediate_23 = usb1_inst_USB_ULPI_DATA_OE_bus[1];
assign intermediate_25 = usb1_inst_USB_ULPI_DATA_OE_bus[2];
assign intermediate_27 = usb1_inst_USB_ULPI_DATA_OE_bus[3];
assign intermediate_29 = usb1_inst_USB_ULPI_DATA_OE_bus[4];
assign intermediate_31 = usb1_inst_USB_ULPI_DATA_OE_bus[5];
assign intermediate_33 = usb1_inst_USB_ULPI_DATA_OE_bus[6];
assign intermediate_35 = usb1_inst_USB_ULPI_DATA_OE_bus[7];

assign intermediate_44 = gpio_inst_GPIO1_PORTA_O_bus[6];
assign intermediate_46 = gpio_inst_GPIO1_PORTA_O_bus[11];
assign intermediate_48 = gpio_inst_GPIO1_PORTA_O_bus[12];
assign intermediate_50 = gpio_inst_GPIO1_PORTA_O_bus[19];
assign intermediate_52 = gpio_inst_GPIO1_PORTA_O_bus[24];
assign intermediate_54 = gpio_inst_GPIO1_PORTA_O_bus[25];

assign intermediate_43 = gpio_inst_GPIO0_PORTA_OE_bus[9];

assign intermediate_56 = gpio_inst_GPIO2_PORTA_O_bus[3];

assign intermediate_42 = gpio_inst_GPIO0_PORTA_O_bus[9];

assign intermediate_57 = gpio_inst_GPIO2_PORTA_OE_bus[3];

assign intermediate_45 = gpio_inst_GPIO1_PORTA_OE_bus[6];
assign intermediate_47 = gpio_inst_GPIO1_PORTA_OE_bus[11];
assign intermediate_49 = gpio_inst_GPIO1_PORTA_OE_bus[12];
assign intermediate_51 = gpio_inst_GPIO1_PORTA_OE_bus[19];
assign intermediate_53 = gpio_inst_GPIO1_PORTA_OE_bus[24];
assign intermediate_55 = gpio_inst_GPIO1_PORTA_OE_bus[25];

assign \gpio_inst~LOANIO0_I0  = gpio_inst_LOANIO0_I_bus[0];
assign \gpio_inst~LOANIO0_I1  = gpio_inst_LOANIO0_I_bus[1];
assign \gpio_inst~LOANIO0_I2  = gpio_inst_LOANIO0_I_bus[2];
assign \gpio_inst~LOANIO0_I3  = gpio_inst_LOANIO0_I_bus[3];
assign \gpio_inst~LOANIO0_I4  = gpio_inst_LOANIO0_I_bus[4];
assign \gpio_inst~LOANIO0_I5  = gpio_inst_LOANIO0_I_bus[5];
assign \gpio_inst~LOANIO0_I6  = gpio_inst_LOANIO0_I_bus[6];
assign \gpio_inst~LOANIO0_I7  = gpio_inst_LOANIO0_I_bus[7];
assign \gpio_inst~LOANIO0_I8  = gpio_inst_LOANIO0_I_bus[8];
assign \gpio_inst~LOANIO0_I9  = gpio_inst_LOANIO0_I_bus[9];
assign \gpio_inst~LOANIO0_I10  = gpio_inst_LOANIO0_I_bus[10];
assign \gpio_inst~LOANIO0_I11  = gpio_inst_LOANIO0_I_bus[11];
assign \gpio_inst~LOANIO0_I12  = gpio_inst_LOANIO0_I_bus[12];
assign \gpio_inst~LOANIO0_I13  = gpio_inst_LOANIO0_I_bus[13];
assign \gpio_inst~LOANIO0_I14  = gpio_inst_LOANIO0_I_bus[14];
assign \gpio_inst~LOANIO0_I15  = gpio_inst_LOANIO0_I_bus[15];
assign \gpio_inst~LOANIO0_I16  = gpio_inst_LOANIO0_I_bus[16];
assign \gpio_inst~LOANIO0_I17  = gpio_inst_LOANIO0_I_bus[17];
assign \gpio_inst~LOANIO0_I18  = gpio_inst_LOANIO0_I_bus[18];
assign \gpio_inst~LOANIO0_I19  = gpio_inst_LOANIO0_I_bus[19];
assign \gpio_inst~LOANIO0_I20  = gpio_inst_LOANIO0_I_bus[20];
assign \gpio_inst~LOANIO0_I21  = gpio_inst_LOANIO0_I_bus[21];
assign \gpio_inst~LOANIO0_I22  = gpio_inst_LOANIO0_I_bus[22];
assign \gpio_inst~LOANIO0_I23  = gpio_inst_LOANIO0_I_bus[23];
assign \gpio_inst~LOANIO0_I24  = gpio_inst_LOANIO0_I_bus[24];
assign \gpio_inst~LOANIO0_I25  = gpio_inst_LOANIO0_I_bus[25];
assign \gpio_inst~LOANIO0_I26  = gpio_inst_LOANIO0_I_bus[26];
assign \gpio_inst~LOANIO0_I27  = gpio_inst_LOANIO0_I_bus[27];
assign \gpio_inst~LOANIO0_I28  = gpio_inst_LOANIO0_I_bus[28];

Computer_System_hps_sdram hps_sdram_inst(
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.GND_port(\~GND~combout ),
	.memory_oct_rzqin(memory_oct_rzqin));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_hps_peripheral_emac emac1_inst(
	.emac_clk_rx(hps_io_emac1_inst_RX_CLK[0]),
	.emac_phy_rxdv(hps_io_emac1_inst_RX_CTL[0]),
	.emac_gmii_mdo_i(hps_io_emac1_inst_MDIO_0),
	.emac_phy_rxd({hps_io_emac1_inst_RXD3[0],hps_io_emac1_inst_RXD2[0],hps_io_emac1_inst_RXD1[0],hps_io_emac1_inst_RXD0[0]}),
	.emac_clk_tx(hps_io_emac1_inst_TX_CLK[0]),
	.emac_phy_tx_oe(hps_io_emac1_inst_TX_CTL[0]),
	.emac_gmii_mdo_o(intermediate_0),
	.emac_gmii_mdo_oe(intermediate_1),
	.emac_gmii_mdc(hps_io_emac1_inst_MDC[0]),
	.emac_phy_txd(emac1_inst_EMAC_PHY_TXD_bus));
defparam emac1_inst.dummy_param = 256;

cyclonev_hps_peripheral_qspi qspi_inst(
	.qspi_mi0(hps_io_qspi_inst_IO0_0),
	.qspi_mi1(hps_io_qspi_inst_IO1_0),
	.qspi_mi2(hps_io_qspi_inst_IO2_0),
	.qspi_mi3(hps_io_qspi_inst_IO3_0),
	.qspi_sclk(hps_io_qspi_inst_CLK[0]),
	.qspi_mo0(intermediate_2),
	.qspi_mo1(intermediate_4),
	.qspi_mo2(intermediate_6),
	.qspi_mo3(intermediate_8),
	.qspi_mo_en_n(qspi_inst_QSPI_MO_EN_N_bus),
	.qspi_ss_n(qspi_inst_QSPI_SS_N_bus));
defparam qspi_inst.dummy_param = 256;

cyclonev_hps_peripheral_sdmmc sdio_inst(
	.sdmmc_fb_clk(gnd),
	.sdmmc_cmd_i(hps_io_sdio_inst_CMD_0),
	.sdmmc_data_i({gnd,gnd,gnd,gnd,hps_io_sdio_inst_D3_0,hps_io_sdio_inst_D2_0,hps_io_sdio_inst_D1_0,hps_io_sdio_inst_D0_0}),
	.sdmmc_pwr_en(\sdio_inst~O_SDMMC_PWR_EN ),
	.sdmmc_cclk(hps_io_sdio_inst_CLK[0]),
	.sdmmc_cmd_o(intermediate_10),
	.sdmmc_cmd_oe(intermediate_11),
	.sdmmc_data_o(sdio_inst_SDMMC_DATA_O_bus),
	.sdmmc_data_oe(sdio_inst_SDMMC_DATA_OE_bus));
defparam sdio_inst.dummy_param = 256;

cyclonev_hps_peripheral_usb usb1_inst(
	.usb_ulpi_clk(hps_io_usb1_inst_CLK[0]),
	.usb_ulpi_dir(hps_io_usb1_inst_DIR[0]),
	.usb_ulpi_nxt(hps_io_usb1_inst_NXT[0]),
	.usb_ulpi_data_i({hps_io_usb1_inst_D7_0,hps_io_usb1_inst_D6_0,hps_io_usb1_inst_D5_0,hps_io_usb1_inst_D4_0,hps_io_usb1_inst_D3_0,hps_io_usb1_inst_D2_0,hps_io_usb1_inst_D1_0,hps_io_usb1_inst_D0_0}),
	.usb_ulpi_stp(hps_io_usb1_inst_STP[0]),
	.usb_ulpi_data_o(usb1_inst_USB_ULPI_DATA_O_bus),
	.usb_ulpi_data_oe(usb1_inst_USB_ULPI_DATA_OE_bus));
defparam usb1_inst.dummy_param = 256;

cyclonev_hps_peripheral_spi_master spim1_inst(
	.spi_master_rxd(hps_io_spim1_inst_MISO[0]),
	.spi_master_sclk(hps_io_spim1_inst_CLK[0]),
	.spi_master_ss_0_n(hps_io_spim1_inst_SS0[0]),
	.spi_master_ss_1_n(),
	.spi_master_txd(intermediate_36),
	.spi_master_ssi_oe_n(intermediate_37));
defparam spim1_inst.dummy_param = 256;

cyclonev_hps_peripheral_uart uart0_inst(
	.uart_cts_n(gnd),
	.uart_rxd(hps_io_uart0_inst_RX[0]),
	.uart_rts_n(\uart0_inst~UARTRTSN ),
	.uart_txd(hps_io_uart0_inst_TX[0]));
defparam uart0_inst.dummy_param = 256;

cyclonev_hps_peripheral_i2c i2c0_inst(
	.i2c_clk(hps_io_i2c0_inst_SCL_0),
	.i2c_data(hps_io_i2c0_inst_SDA_0),
	.i2c_clk_oe(intermediate_39),
	.i2c_data_oe(intermediate_38));
defparam i2c0_inst.dummy_param = 256;

cyclonev_hps_peripheral_i2c i2c1_inst(
	.i2c_clk(hps_io_i2c1_inst_SCL_0),
	.i2c_data(hps_io_i2c1_inst_SDA_0),
	.i2c_clk_oe(intermediate_41),
	.i2c_data_oe(intermediate_40));
defparam i2c1_inst.dummy_param = 256;

cyclonev_hps_peripheral_gpio gpio_inst(
	.gpio0_porta_i({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO09_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.gpio1_porta_i({gnd,gnd,gnd,hps_io_gpio_inst_GPIO54_0,hps_io_gpio_inst_GPIO53_0,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO48_0,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO41_0,hps_io_gpio_inst_GPIO40_0,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO35_0,gnd,gnd,gnd,gnd,gnd,gnd}),
	.gpio2_porta_i({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO61_0,gnd,gnd,gnd}),
	.loanio0_o(29'b00000000000000000000000000000),
	.loanio0_oe(29'b00000000000000000000000000000),
	.loanio1_o(29'b00000000000000000000000000000),
	.loanio1_oe(29'b00000000000000000000000000000),
	.loanio2_o(29'b00000000000000000000000000000),
	.loanio2_oe(29'b00000000000000000000000000000),
	.loanio0_i(gpio_inst_LOANIO0_I_bus),
	.loanio1_i(),
	.loanio2_i(),
	.gpio0_porta_o(gpio_inst_GPIO0_PORTA_O_bus),
	.gpio0_porta_oe(gpio_inst_GPIO0_PORTA_OE_bus),
	.gpio1_porta_o(gpio_inst_GPIO1_PORTA_O_bus),
	.gpio1_porta_oe(gpio_inst_GPIO1_PORTA_OE_bus),
	.gpio2_porta_o(gpio_inst_GPIO2_PORTA_O_bus),
	.gpio2_porta_oe(gpio_inst_GPIO2_PORTA_OE_bus));
defparam gpio_inst.dummy_param = 256;

endmodule

module Computer_System_hps_sdram (
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	GND_port,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	GND_port;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pll|afi_clk ;
wire \pll|pll_write_clk ;
wire \p0|umemphy|afi_cal_fail ;
wire \p0|umemphy|afi_cal_success ;
wire \p0|umemphy|afi_rdata_valid[0] ;
wire \p0|umemphy|ctl_reset_n ;
wire \p0|umemphy|afi_rdata[0] ;
wire \p0|umemphy|afi_rdata[1] ;
wire \p0|umemphy|afi_rdata[2] ;
wire \p0|umemphy|afi_rdata[3] ;
wire \p0|umemphy|afi_rdata[4] ;
wire \p0|umemphy|afi_rdata[5] ;
wire \p0|umemphy|afi_rdata[6] ;
wire \p0|umemphy|afi_rdata[7] ;
wire \p0|umemphy|afi_rdata[8] ;
wire \p0|umemphy|afi_rdata[9] ;
wire \p0|umemphy|afi_rdata[10] ;
wire \p0|umemphy|afi_rdata[11] ;
wire \p0|umemphy|afi_rdata[12] ;
wire \p0|umemphy|afi_rdata[13] ;
wire \p0|umemphy|afi_rdata[14] ;
wire \p0|umemphy|afi_rdata[15] ;
wire \p0|umemphy|afi_rdata[16] ;
wire \p0|umemphy|afi_rdata[17] ;
wire \p0|umemphy|afi_rdata[18] ;
wire \p0|umemphy|afi_rdata[19] ;
wire \p0|umemphy|afi_rdata[20] ;
wire \p0|umemphy|afi_rdata[21] ;
wire \p0|umemphy|afi_rdata[22] ;
wire \p0|umemphy|afi_rdata[23] ;
wire \p0|umemphy|afi_rdata[24] ;
wire \p0|umemphy|afi_rdata[25] ;
wire \p0|umemphy|afi_rdata[26] ;
wire \p0|umemphy|afi_rdata[27] ;
wire \p0|umemphy|afi_rdata[28] ;
wire \p0|umemphy|afi_rdata[29] ;
wire \p0|umemphy|afi_rdata[30] ;
wire \p0|umemphy|afi_rdata[31] ;
wire \p0|umemphy|afi_rdata[32] ;
wire \p0|umemphy|afi_rdata[33] ;
wire \p0|umemphy|afi_rdata[34] ;
wire \p0|umemphy|afi_rdata[35] ;
wire \p0|umemphy|afi_rdata[36] ;
wire \p0|umemphy|afi_rdata[37] ;
wire \p0|umemphy|afi_rdata[38] ;
wire \p0|umemphy|afi_rdata[39] ;
wire \p0|umemphy|afi_rdata[40] ;
wire \p0|umemphy|afi_rdata[41] ;
wire \p0|umemphy|afi_rdata[42] ;
wire \p0|umemphy|afi_rdata[43] ;
wire \p0|umemphy|afi_rdata[44] ;
wire \p0|umemphy|afi_rdata[45] ;
wire \p0|umemphy|afi_rdata[46] ;
wire \p0|umemphy|afi_rdata[47] ;
wire \p0|umemphy|afi_rdata[48] ;
wire \p0|umemphy|afi_rdata[49] ;
wire \p0|umemphy|afi_rdata[50] ;
wire \p0|umemphy|afi_rdata[51] ;
wire \p0|umemphy|afi_rdata[52] ;
wire \p0|umemphy|afi_rdata[53] ;
wire \p0|umemphy|afi_rdata[54] ;
wire \p0|umemphy|afi_rdata[55] ;
wire \p0|umemphy|afi_rdata[56] ;
wire \p0|umemphy|afi_rdata[57] ;
wire \p0|umemphy|afi_rdata[58] ;
wire \p0|umemphy|afi_rdata[59] ;
wire \p0|umemphy|afi_rdata[60] ;
wire \p0|umemphy|afi_rdata[61] ;
wire \p0|umemphy|afi_rdata[62] ;
wire \p0|umemphy|afi_rdata[63] ;
wire \p0|umemphy|afi_rdata[64] ;
wire \p0|umemphy|afi_rdata[65] ;
wire \p0|umemphy|afi_rdata[66] ;
wire \p0|umemphy|afi_rdata[67] ;
wire \p0|umemphy|afi_rdata[68] ;
wire \p0|umemphy|afi_rdata[69] ;
wire \p0|umemphy|afi_rdata[70] ;
wire \p0|umemphy|afi_rdata[71] ;
wire \p0|umemphy|afi_rdata[72] ;
wire \p0|umemphy|afi_rdata[73] ;
wire \p0|umemphy|afi_rdata[74] ;
wire \p0|umemphy|afi_rdata[75] ;
wire \p0|umemphy|afi_rdata[76] ;
wire \p0|umemphy|afi_rdata[77] ;
wire \p0|umemphy|afi_rdata[78] ;
wire \p0|umemphy|afi_rdata[79] ;
wire \p0|umemphy|afi_wlat[0] ;
wire \p0|umemphy|afi_wlat[1] ;
wire \p0|umemphy|afi_wlat[2] ;
wire \p0|umemphy|afi_wlat[3] ;
wire \c0|afi_cas_n[0] ;
wire \c0|afi_ras_n[0] ;
wire \c0|afi_rst_n[0] ;
wire \c0|afi_we_n[0] ;
wire \c0|afi_addr[0] ;
wire \c0|afi_addr[1] ;
wire \c0|afi_addr[2] ;
wire \c0|afi_addr[3] ;
wire \c0|afi_addr[4] ;
wire \c0|afi_addr[5] ;
wire \c0|afi_addr[6] ;
wire \c0|afi_addr[7] ;
wire \c0|afi_addr[8] ;
wire \c0|afi_addr[9] ;
wire \c0|afi_addr[10] ;
wire \c0|afi_addr[11] ;
wire \c0|afi_addr[12] ;
wire \c0|afi_addr[13] ;
wire \c0|afi_addr[14] ;
wire \c0|afi_addr[15] ;
wire \c0|afi_addr[16] ;
wire \c0|afi_addr[17] ;
wire \c0|afi_addr[18] ;
wire \c0|afi_addr[19] ;
wire \c0|afi_ba[0] ;
wire \c0|afi_ba[1] ;
wire \c0|afi_ba[2] ;
wire \c0|afi_cke[0] ;
wire \c0|afi_cke[1] ;
wire \c0|afi_cs_n[0] ;
wire \c0|afi_cs_n[1] ;
wire \c0|afi_dm_int[0] ;
wire \c0|afi_dm_int[1] ;
wire \c0|afi_dm_int[2] ;
wire \c0|afi_dm_int[3] ;
wire \c0|afi_dm_int[4] ;
wire \c0|afi_dm_int[5] ;
wire \c0|afi_dm_int[6] ;
wire \c0|afi_dm_int[7] ;
wire \c0|afi_dm_int[8] ;
wire \c0|afi_dm_int[9] ;
wire \c0|afi_dqs_burst[0] ;
wire \c0|afi_dqs_burst[1] ;
wire \c0|afi_dqs_burst[2] ;
wire \c0|afi_dqs_burst[3] ;
wire \c0|afi_dqs_burst[4] ;
wire \c0|afi_odt[0] ;
wire \c0|afi_odt[1] ;
wire \c0|afi_rdata_en[0] ;
wire \c0|afi_rdata_en[1] ;
wire \c0|afi_rdata_en[2] ;
wire \c0|afi_rdata_en[3] ;
wire \c0|afi_rdata_en[4] ;
wire \c0|afi_rdata_en_full[0] ;
wire \c0|afi_rdata_en_full[1] ;
wire \c0|afi_rdata_en_full[2] ;
wire \c0|afi_rdata_en_full[3] ;
wire \c0|afi_rdata_en_full[4] ;
wire \c0|afi_wdata_int[0] ;
wire \c0|afi_wdata_int[1] ;
wire \c0|afi_wdata_int[2] ;
wire \c0|afi_wdata_int[3] ;
wire \c0|afi_wdata_int[4] ;
wire \c0|afi_wdata_int[5] ;
wire \c0|afi_wdata_int[6] ;
wire \c0|afi_wdata_int[7] ;
wire \c0|afi_wdata_int[8] ;
wire \c0|afi_wdata_int[9] ;
wire \c0|afi_wdata_int[10] ;
wire \c0|afi_wdata_int[11] ;
wire \c0|afi_wdata_int[12] ;
wire \c0|afi_wdata_int[13] ;
wire \c0|afi_wdata_int[14] ;
wire \c0|afi_wdata_int[15] ;
wire \c0|afi_wdata_int[16] ;
wire \c0|afi_wdata_int[17] ;
wire \c0|afi_wdata_int[18] ;
wire \c0|afi_wdata_int[19] ;
wire \c0|afi_wdata_int[20] ;
wire \c0|afi_wdata_int[21] ;
wire \c0|afi_wdata_int[22] ;
wire \c0|afi_wdata_int[23] ;
wire \c0|afi_wdata_int[24] ;
wire \c0|afi_wdata_int[25] ;
wire \c0|afi_wdata_int[26] ;
wire \c0|afi_wdata_int[27] ;
wire \c0|afi_wdata_int[28] ;
wire \c0|afi_wdata_int[29] ;
wire \c0|afi_wdata_int[30] ;
wire \c0|afi_wdata_int[31] ;
wire \c0|afi_wdata_int[32] ;
wire \c0|afi_wdata_int[33] ;
wire \c0|afi_wdata_int[34] ;
wire \c0|afi_wdata_int[35] ;
wire \c0|afi_wdata_int[36] ;
wire \c0|afi_wdata_int[37] ;
wire \c0|afi_wdata_int[38] ;
wire \c0|afi_wdata_int[39] ;
wire \c0|afi_wdata_int[40] ;
wire \c0|afi_wdata_int[41] ;
wire \c0|afi_wdata_int[42] ;
wire \c0|afi_wdata_int[43] ;
wire \c0|afi_wdata_int[44] ;
wire \c0|afi_wdata_int[45] ;
wire \c0|afi_wdata_int[46] ;
wire \c0|afi_wdata_int[47] ;
wire \c0|afi_wdata_int[48] ;
wire \c0|afi_wdata_int[49] ;
wire \c0|afi_wdata_int[50] ;
wire \c0|afi_wdata_int[51] ;
wire \c0|afi_wdata_int[52] ;
wire \c0|afi_wdata_int[53] ;
wire \c0|afi_wdata_int[54] ;
wire \c0|afi_wdata_int[55] ;
wire \c0|afi_wdata_int[56] ;
wire \c0|afi_wdata_int[57] ;
wire \c0|afi_wdata_int[58] ;
wire \c0|afi_wdata_int[59] ;
wire \c0|afi_wdata_int[60] ;
wire \c0|afi_wdata_int[61] ;
wire \c0|afi_wdata_int[62] ;
wire \c0|afi_wdata_int[63] ;
wire \c0|afi_wdata_int[64] ;
wire \c0|afi_wdata_int[65] ;
wire \c0|afi_wdata_int[66] ;
wire \c0|afi_wdata_int[67] ;
wire \c0|afi_wdata_int[68] ;
wire \c0|afi_wdata_int[69] ;
wire \c0|afi_wdata_int[70] ;
wire \c0|afi_wdata_int[71] ;
wire \c0|afi_wdata_int[72] ;
wire \c0|afi_wdata_int[73] ;
wire \c0|afi_wdata_int[74] ;
wire \c0|afi_wdata_int[75] ;
wire \c0|afi_wdata_int[76] ;
wire \c0|afi_wdata_int[77] ;
wire \c0|afi_wdata_int[78] ;
wire \c0|afi_wdata_int[79] ;
wire \c0|afi_wdata_valid[0] ;
wire \c0|afi_wdata_valid[1] ;
wire \c0|afi_wdata_valid[2] ;
wire \c0|afi_wdata_valid[3] ;
wire \c0|afi_wdata_valid[4] ;
wire \c0|cfg_addlat_wire[0] ;
wire \c0|cfg_addlat_wire[1] ;
wire \c0|cfg_addlat_wire[2] ;
wire \c0|cfg_addlat_wire[3] ;
wire \c0|cfg_addlat_wire[4] ;
wire \c0|cfg_bankaddrwidth_wire[0] ;
wire \c0|cfg_bankaddrwidth_wire[1] ;
wire \c0|cfg_bankaddrwidth_wire[2] ;
wire \c0|cfg_caswrlat_wire[0] ;
wire \c0|cfg_caswrlat_wire[1] ;
wire \c0|cfg_caswrlat_wire[2] ;
wire \c0|cfg_caswrlat_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[0] ;
wire \c0|cfg_coladdrwidth_wire[1] ;
wire \c0|cfg_coladdrwidth_wire[2] ;
wire \c0|cfg_coladdrwidth_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[4] ;
wire \c0|cfg_csaddrwidth_wire[0] ;
wire \c0|cfg_csaddrwidth_wire[1] ;
wire \c0|cfg_csaddrwidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[0] ;
wire \c0|cfg_devicewidth_wire[1] ;
wire \c0|cfg_devicewidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[0] ;
wire \c0|cfg_interfacewidth_wire[1] ;
wire \c0|cfg_interfacewidth_wire[2] ;
wire \c0|cfg_interfacewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[4] ;
wire \c0|cfg_interfacewidth_wire[5] ;
wire \c0|cfg_interfacewidth_wire[6] ;
wire \c0|cfg_interfacewidth_wire[7] ;
wire \c0|cfg_rowaddrwidth_wire[0] ;
wire \c0|cfg_rowaddrwidth_wire[1] ;
wire \c0|cfg_rowaddrwidth_wire[2] ;
wire \c0|cfg_rowaddrwidth_wire[3] ;
wire \c0|cfg_rowaddrwidth_wire[4] ;
wire \c0|cfg_tcl_wire[0] ;
wire \c0|cfg_tcl_wire[1] ;
wire \c0|cfg_tcl_wire[2] ;
wire \c0|cfg_tcl_wire[3] ;
wire \c0|cfg_tcl_wire[4] ;
wire \c0|cfg_tmrd_wire[0] ;
wire \c0|cfg_tmrd_wire[1] ;
wire \c0|cfg_tmrd_wire[2] ;
wire \c0|cfg_tmrd_wire[3] ;
wire \c0|cfg_trefi_wire[0] ;
wire \c0|cfg_trefi_wire[1] ;
wire \c0|cfg_trefi_wire[2] ;
wire \c0|cfg_trefi_wire[3] ;
wire \c0|cfg_trefi_wire[4] ;
wire \c0|cfg_trefi_wire[5] ;
wire \c0|cfg_trefi_wire[6] ;
wire \c0|cfg_trefi_wire[7] ;
wire \c0|cfg_trefi_wire[8] ;
wire \c0|cfg_trefi_wire[9] ;
wire \c0|cfg_trefi_wire[10] ;
wire \c0|cfg_trefi_wire[11] ;
wire \c0|cfg_trefi_wire[12] ;
wire \c0|cfg_trfc_wire[0] ;
wire \c0|cfg_trfc_wire[1] ;
wire \c0|cfg_trfc_wire[2] ;
wire \c0|cfg_trfc_wire[3] ;
wire \c0|cfg_trfc_wire[4] ;
wire \c0|cfg_trfc_wire[5] ;
wire \c0|cfg_trfc_wire[6] ;
wire \c0|cfg_trfc_wire[7] ;
wire \c0|cfg_twr_wire[0] ;
wire \c0|cfg_twr_wire[1] ;
wire \c0|cfg_twr_wire[2] ;
wire \c0|cfg_twr_wire[3] ;
wire \c0|afi_mem_clk_disable[0] ;
wire \c0|cfg_dramconfig_wire[0] ;
wire \c0|cfg_dramconfig_wire[1] ;
wire \c0|cfg_dramconfig_wire[2] ;
wire \c0|cfg_dramconfig_wire[3] ;
wire \c0|cfg_dramconfig_wire[4] ;
wire \c0|cfg_dramconfig_wire[5] ;
wire \c0|cfg_dramconfig_wire[6] ;
wire \c0|cfg_dramconfig_wire[7] ;
wire \c0|cfg_dramconfig_wire[8] ;
wire \c0|cfg_dramconfig_wire[9] ;
wire \c0|cfg_dramconfig_wire[10] ;
wire \c0|cfg_dramconfig_wire[11] ;
wire \c0|cfg_dramconfig_wire[12] ;
wire \c0|cfg_dramconfig_wire[13] ;
wire \c0|cfg_dramconfig_wire[14] ;
wire \c0|cfg_dramconfig_wire[15] ;
wire \c0|cfg_dramconfig_wire[16] ;
wire \c0|cfg_dramconfig_wire[17] ;
wire \c0|cfg_dramconfig_wire[18] ;
wire \c0|cfg_dramconfig_wire[19] ;
wire \c0|cfg_dramconfig_wire[20] ;
wire \p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ;
wire \dll|dll_delayctrl[0] ;
wire \dll|dll_delayctrl[1] ;
wire \dll|dll_delayctrl[2] ;
wire \dll|dll_delayctrl[3] ;
wire \dll|dll_delayctrl[4] ;
wire \dll|dll_delayctrl[5] ;
wire \dll|dll_delayctrl[6] ;


Computer_System_hps_sdram_p0 p0(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid_0(\p0|umemphy|afi_rdata_valid[0] ),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata_0(\p0|umemphy|afi_rdata[0] ),
	.afi_rdata_1(\p0|umemphy|afi_rdata[1] ),
	.afi_rdata_2(\p0|umemphy|afi_rdata[2] ),
	.afi_rdata_3(\p0|umemphy|afi_rdata[3] ),
	.afi_rdata_4(\p0|umemphy|afi_rdata[4] ),
	.afi_rdata_5(\p0|umemphy|afi_rdata[5] ),
	.afi_rdata_6(\p0|umemphy|afi_rdata[6] ),
	.afi_rdata_7(\p0|umemphy|afi_rdata[7] ),
	.afi_rdata_8(\p0|umemphy|afi_rdata[8] ),
	.afi_rdata_9(\p0|umemphy|afi_rdata[9] ),
	.afi_rdata_10(\p0|umemphy|afi_rdata[10] ),
	.afi_rdata_11(\p0|umemphy|afi_rdata[11] ),
	.afi_rdata_12(\p0|umemphy|afi_rdata[12] ),
	.afi_rdata_13(\p0|umemphy|afi_rdata[13] ),
	.afi_rdata_14(\p0|umemphy|afi_rdata[14] ),
	.afi_rdata_15(\p0|umemphy|afi_rdata[15] ),
	.afi_rdata_16(\p0|umemphy|afi_rdata[16] ),
	.afi_rdata_17(\p0|umemphy|afi_rdata[17] ),
	.afi_rdata_18(\p0|umemphy|afi_rdata[18] ),
	.afi_rdata_19(\p0|umemphy|afi_rdata[19] ),
	.afi_rdata_20(\p0|umemphy|afi_rdata[20] ),
	.afi_rdata_21(\p0|umemphy|afi_rdata[21] ),
	.afi_rdata_22(\p0|umemphy|afi_rdata[22] ),
	.afi_rdata_23(\p0|umemphy|afi_rdata[23] ),
	.afi_rdata_24(\p0|umemphy|afi_rdata[24] ),
	.afi_rdata_25(\p0|umemphy|afi_rdata[25] ),
	.afi_rdata_26(\p0|umemphy|afi_rdata[26] ),
	.afi_rdata_27(\p0|umemphy|afi_rdata[27] ),
	.afi_rdata_28(\p0|umemphy|afi_rdata[28] ),
	.afi_rdata_29(\p0|umemphy|afi_rdata[29] ),
	.afi_rdata_30(\p0|umemphy|afi_rdata[30] ),
	.afi_rdata_31(\p0|umemphy|afi_rdata[31] ),
	.afi_rdata_32(\p0|umemphy|afi_rdata[32] ),
	.afi_rdata_33(\p0|umemphy|afi_rdata[33] ),
	.afi_rdata_34(\p0|umemphy|afi_rdata[34] ),
	.afi_rdata_35(\p0|umemphy|afi_rdata[35] ),
	.afi_rdata_36(\p0|umemphy|afi_rdata[36] ),
	.afi_rdata_37(\p0|umemphy|afi_rdata[37] ),
	.afi_rdata_38(\p0|umemphy|afi_rdata[38] ),
	.afi_rdata_39(\p0|umemphy|afi_rdata[39] ),
	.afi_rdata_40(\p0|umemphy|afi_rdata[40] ),
	.afi_rdata_41(\p0|umemphy|afi_rdata[41] ),
	.afi_rdata_42(\p0|umemphy|afi_rdata[42] ),
	.afi_rdata_43(\p0|umemphy|afi_rdata[43] ),
	.afi_rdata_44(\p0|umemphy|afi_rdata[44] ),
	.afi_rdata_45(\p0|umemphy|afi_rdata[45] ),
	.afi_rdata_46(\p0|umemphy|afi_rdata[46] ),
	.afi_rdata_47(\p0|umemphy|afi_rdata[47] ),
	.afi_rdata_48(\p0|umemphy|afi_rdata[48] ),
	.afi_rdata_49(\p0|umemphy|afi_rdata[49] ),
	.afi_rdata_50(\p0|umemphy|afi_rdata[50] ),
	.afi_rdata_51(\p0|umemphy|afi_rdata[51] ),
	.afi_rdata_52(\p0|umemphy|afi_rdata[52] ),
	.afi_rdata_53(\p0|umemphy|afi_rdata[53] ),
	.afi_rdata_54(\p0|umemphy|afi_rdata[54] ),
	.afi_rdata_55(\p0|umemphy|afi_rdata[55] ),
	.afi_rdata_56(\p0|umemphy|afi_rdata[56] ),
	.afi_rdata_57(\p0|umemphy|afi_rdata[57] ),
	.afi_rdata_58(\p0|umemphy|afi_rdata[58] ),
	.afi_rdata_59(\p0|umemphy|afi_rdata[59] ),
	.afi_rdata_60(\p0|umemphy|afi_rdata[60] ),
	.afi_rdata_61(\p0|umemphy|afi_rdata[61] ),
	.afi_rdata_62(\p0|umemphy|afi_rdata[62] ),
	.afi_rdata_63(\p0|umemphy|afi_rdata[63] ),
	.afi_rdata_64(\p0|umemphy|afi_rdata[64] ),
	.afi_rdata_65(\p0|umemphy|afi_rdata[65] ),
	.afi_rdata_66(\p0|umemphy|afi_rdata[66] ),
	.afi_rdata_67(\p0|umemphy|afi_rdata[67] ),
	.afi_rdata_68(\p0|umemphy|afi_rdata[68] ),
	.afi_rdata_69(\p0|umemphy|afi_rdata[69] ),
	.afi_rdata_70(\p0|umemphy|afi_rdata[70] ),
	.afi_rdata_71(\p0|umemphy|afi_rdata[71] ),
	.afi_rdata_72(\p0|umemphy|afi_rdata[72] ),
	.afi_rdata_73(\p0|umemphy|afi_rdata[73] ),
	.afi_rdata_74(\p0|umemphy|afi_rdata[74] ),
	.afi_rdata_75(\p0|umemphy|afi_rdata[75] ),
	.afi_rdata_76(\p0|umemphy|afi_rdata[76] ),
	.afi_rdata_77(\p0|umemphy|afi_rdata[77] ),
	.afi_rdata_78(\p0|umemphy|afi_rdata[78] ),
	.afi_rdata_79(\p0|umemphy|afi_rdata[79] ),
	.afi_wlat_0(\p0|umemphy|afi_wlat[0] ),
	.afi_wlat_1(\p0|umemphy|afi_wlat[1] ),
	.afi_wlat_2(\p0|umemphy|afi_wlat[2] ),
	.afi_wlat_3(\p0|umemphy|afi_wlat[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n_0(\c0|afi_cas_n[0] ),
	.afi_ras_n_0(\c0|afi_ras_n[0] ),
	.afi_rst_n_0(\c0|afi_rst_n[0] ),
	.afi_we_n_0(\c0|afi_we_n[0] ),
	.afi_addr_0(\c0|afi_addr[0] ),
	.afi_addr_1(\c0|afi_addr[1] ),
	.afi_addr_2(\c0|afi_addr[2] ),
	.afi_addr_3(\c0|afi_addr[3] ),
	.afi_addr_4(\c0|afi_addr[4] ),
	.afi_addr_5(\c0|afi_addr[5] ),
	.afi_addr_6(\c0|afi_addr[6] ),
	.afi_addr_7(\c0|afi_addr[7] ),
	.afi_addr_8(\c0|afi_addr[8] ),
	.afi_addr_9(\c0|afi_addr[9] ),
	.afi_addr_10(\c0|afi_addr[10] ),
	.afi_addr_11(\c0|afi_addr[11] ),
	.afi_addr_12(\c0|afi_addr[12] ),
	.afi_addr_13(\c0|afi_addr[13] ),
	.afi_addr_14(\c0|afi_addr[14] ),
	.afi_addr_15(\c0|afi_addr[15] ),
	.afi_addr_16(\c0|afi_addr[16] ),
	.afi_addr_17(\c0|afi_addr[17] ),
	.afi_addr_18(\c0|afi_addr[18] ),
	.afi_addr_19(\c0|afi_addr[19] ),
	.afi_ba_0(\c0|afi_ba[0] ),
	.afi_ba_1(\c0|afi_ba[1] ),
	.afi_ba_2(\c0|afi_ba[2] ),
	.afi_cke_0(\c0|afi_cke[0] ),
	.afi_cke_1(\c0|afi_cke[1] ),
	.afi_cs_n_0(\c0|afi_cs_n[0] ),
	.afi_cs_n_1(\c0|afi_cs_n[1] ),
	.afi_dm_int_0(\c0|afi_dm_int[0] ),
	.afi_dm_int_1(\c0|afi_dm_int[1] ),
	.afi_dm_int_2(\c0|afi_dm_int[2] ),
	.afi_dm_int_3(\c0|afi_dm_int[3] ),
	.afi_dm_int_4(\c0|afi_dm_int[4] ),
	.afi_dm_int_5(\c0|afi_dm_int[5] ),
	.afi_dm_int_6(\c0|afi_dm_int[6] ),
	.afi_dm_int_7(\c0|afi_dm_int[7] ),
	.afi_dm_int_8(\c0|afi_dm_int[8] ),
	.afi_dm_int_9(\c0|afi_dm_int[9] ),
	.afi_dqs_burst_0(\c0|afi_dqs_burst[0] ),
	.afi_dqs_burst_1(\c0|afi_dqs_burst[1] ),
	.afi_dqs_burst_2(\c0|afi_dqs_burst[2] ),
	.afi_dqs_burst_3(\c0|afi_dqs_burst[3] ),
	.afi_dqs_burst_4(\c0|afi_dqs_burst[4] ),
	.afi_odt_0(\c0|afi_odt[0] ),
	.afi_odt_1(\c0|afi_odt[1] ),
	.afi_rdata_en_0(\c0|afi_rdata_en[0] ),
	.afi_rdata_en_1(\c0|afi_rdata_en[1] ),
	.afi_rdata_en_2(\c0|afi_rdata_en[2] ),
	.afi_rdata_en_3(\c0|afi_rdata_en[3] ),
	.afi_rdata_en_4(\c0|afi_rdata_en[4] ),
	.afi_rdata_en_full_0(\c0|afi_rdata_en_full[0] ),
	.afi_rdata_en_full_1(\c0|afi_rdata_en_full[1] ),
	.afi_rdata_en_full_2(\c0|afi_rdata_en_full[2] ),
	.afi_rdata_en_full_3(\c0|afi_rdata_en_full[3] ),
	.afi_rdata_en_full_4(\c0|afi_rdata_en_full[4] ),
	.afi_wdata_int_0(\c0|afi_wdata_int[0] ),
	.afi_wdata_int_1(\c0|afi_wdata_int[1] ),
	.afi_wdata_int_2(\c0|afi_wdata_int[2] ),
	.afi_wdata_int_3(\c0|afi_wdata_int[3] ),
	.afi_wdata_int_4(\c0|afi_wdata_int[4] ),
	.afi_wdata_int_5(\c0|afi_wdata_int[5] ),
	.afi_wdata_int_6(\c0|afi_wdata_int[6] ),
	.afi_wdata_int_7(\c0|afi_wdata_int[7] ),
	.afi_wdata_int_8(\c0|afi_wdata_int[8] ),
	.afi_wdata_int_9(\c0|afi_wdata_int[9] ),
	.afi_wdata_int_10(\c0|afi_wdata_int[10] ),
	.afi_wdata_int_11(\c0|afi_wdata_int[11] ),
	.afi_wdata_int_12(\c0|afi_wdata_int[12] ),
	.afi_wdata_int_13(\c0|afi_wdata_int[13] ),
	.afi_wdata_int_14(\c0|afi_wdata_int[14] ),
	.afi_wdata_int_15(\c0|afi_wdata_int[15] ),
	.afi_wdata_int_16(\c0|afi_wdata_int[16] ),
	.afi_wdata_int_17(\c0|afi_wdata_int[17] ),
	.afi_wdata_int_18(\c0|afi_wdata_int[18] ),
	.afi_wdata_int_19(\c0|afi_wdata_int[19] ),
	.afi_wdata_int_20(\c0|afi_wdata_int[20] ),
	.afi_wdata_int_21(\c0|afi_wdata_int[21] ),
	.afi_wdata_int_22(\c0|afi_wdata_int[22] ),
	.afi_wdata_int_23(\c0|afi_wdata_int[23] ),
	.afi_wdata_int_24(\c0|afi_wdata_int[24] ),
	.afi_wdata_int_25(\c0|afi_wdata_int[25] ),
	.afi_wdata_int_26(\c0|afi_wdata_int[26] ),
	.afi_wdata_int_27(\c0|afi_wdata_int[27] ),
	.afi_wdata_int_28(\c0|afi_wdata_int[28] ),
	.afi_wdata_int_29(\c0|afi_wdata_int[29] ),
	.afi_wdata_int_30(\c0|afi_wdata_int[30] ),
	.afi_wdata_int_31(\c0|afi_wdata_int[31] ),
	.afi_wdata_int_32(\c0|afi_wdata_int[32] ),
	.afi_wdata_int_33(\c0|afi_wdata_int[33] ),
	.afi_wdata_int_34(\c0|afi_wdata_int[34] ),
	.afi_wdata_int_35(\c0|afi_wdata_int[35] ),
	.afi_wdata_int_36(\c0|afi_wdata_int[36] ),
	.afi_wdata_int_37(\c0|afi_wdata_int[37] ),
	.afi_wdata_int_38(\c0|afi_wdata_int[38] ),
	.afi_wdata_int_39(\c0|afi_wdata_int[39] ),
	.afi_wdata_int_40(\c0|afi_wdata_int[40] ),
	.afi_wdata_int_41(\c0|afi_wdata_int[41] ),
	.afi_wdata_int_42(\c0|afi_wdata_int[42] ),
	.afi_wdata_int_43(\c0|afi_wdata_int[43] ),
	.afi_wdata_int_44(\c0|afi_wdata_int[44] ),
	.afi_wdata_int_45(\c0|afi_wdata_int[45] ),
	.afi_wdata_int_46(\c0|afi_wdata_int[46] ),
	.afi_wdata_int_47(\c0|afi_wdata_int[47] ),
	.afi_wdata_int_48(\c0|afi_wdata_int[48] ),
	.afi_wdata_int_49(\c0|afi_wdata_int[49] ),
	.afi_wdata_int_50(\c0|afi_wdata_int[50] ),
	.afi_wdata_int_51(\c0|afi_wdata_int[51] ),
	.afi_wdata_int_52(\c0|afi_wdata_int[52] ),
	.afi_wdata_int_53(\c0|afi_wdata_int[53] ),
	.afi_wdata_int_54(\c0|afi_wdata_int[54] ),
	.afi_wdata_int_55(\c0|afi_wdata_int[55] ),
	.afi_wdata_int_56(\c0|afi_wdata_int[56] ),
	.afi_wdata_int_57(\c0|afi_wdata_int[57] ),
	.afi_wdata_int_58(\c0|afi_wdata_int[58] ),
	.afi_wdata_int_59(\c0|afi_wdata_int[59] ),
	.afi_wdata_int_60(\c0|afi_wdata_int[60] ),
	.afi_wdata_int_61(\c0|afi_wdata_int[61] ),
	.afi_wdata_int_62(\c0|afi_wdata_int[62] ),
	.afi_wdata_int_63(\c0|afi_wdata_int[63] ),
	.afi_wdata_int_64(\c0|afi_wdata_int[64] ),
	.afi_wdata_int_65(\c0|afi_wdata_int[65] ),
	.afi_wdata_int_66(\c0|afi_wdata_int[66] ),
	.afi_wdata_int_67(\c0|afi_wdata_int[67] ),
	.afi_wdata_int_68(\c0|afi_wdata_int[68] ),
	.afi_wdata_int_69(\c0|afi_wdata_int[69] ),
	.afi_wdata_int_70(\c0|afi_wdata_int[70] ),
	.afi_wdata_int_71(\c0|afi_wdata_int[71] ),
	.afi_wdata_int_72(\c0|afi_wdata_int[72] ),
	.afi_wdata_int_73(\c0|afi_wdata_int[73] ),
	.afi_wdata_int_74(\c0|afi_wdata_int[74] ),
	.afi_wdata_int_75(\c0|afi_wdata_int[75] ),
	.afi_wdata_int_76(\c0|afi_wdata_int[76] ),
	.afi_wdata_int_77(\c0|afi_wdata_int[77] ),
	.afi_wdata_int_78(\c0|afi_wdata_int[78] ),
	.afi_wdata_int_79(\c0|afi_wdata_int[79] ),
	.afi_wdata_valid_0(\c0|afi_wdata_valid[0] ),
	.afi_wdata_valid_1(\c0|afi_wdata_valid[1] ),
	.afi_wdata_valid_2(\c0|afi_wdata_valid[2] ),
	.afi_wdata_valid_3(\c0|afi_wdata_valid[3] ),
	.afi_wdata_valid_4(\c0|afi_wdata_valid[4] ),
	.cfg_addlat_wire_0(\c0|cfg_addlat_wire[0] ),
	.cfg_addlat_wire_1(\c0|cfg_addlat_wire[1] ),
	.cfg_addlat_wire_2(\c0|cfg_addlat_wire[2] ),
	.cfg_addlat_wire_3(\c0|cfg_addlat_wire[3] ),
	.cfg_addlat_wire_4(\c0|cfg_addlat_wire[4] ),
	.cfg_bankaddrwidth_wire_0(\c0|cfg_bankaddrwidth_wire[0] ),
	.cfg_bankaddrwidth_wire_1(\c0|cfg_bankaddrwidth_wire[1] ),
	.cfg_bankaddrwidth_wire_2(\c0|cfg_bankaddrwidth_wire[2] ),
	.cfg_caswrlat_wire_0(\c0|cfg_caswrlat_wire[0] ),
	.cfg_caswrlat_wire_1(\c0|cfg_caswrlat_wire[1] ),
	.cfg_caswrlat_wire_2(\c0|cfg_caswrlat_wire[2] ),
	.cfg_caswrlat_wire_3(\c0|cfg_caswrlat_wire[3] ),
	.cfg_coladdrwidth_wire_0(\c0|cfg_coladdrwidth_wire[0] ),
	.cfg_coladdrwidth_wire_1(\c0|cfg_coladdrwidth_wire[1] ),
	.cfg_coladdrwidth_wire_2(\c0|cfg_coladdrwidth_wire[2] ),
	.cfg_coladdrwidth_wire_3(\c0|cfg_coladdrwidth_wire[3] ),
	.cfg_coladdrwidth_wire_4(\c0|cfg_coladdrwidth_wire[4] ),
	.cfg_csaddrwidth_wire_0(\c0|cfg_csaddrwidth_wire[0] ),
	.cfg_csaddrwidth_wire_1(\c0|cfg_csaddrwidth_wire[1] ),
	.cfg_csaddrwidth_wire_2(\c0|cfg_csaddrwidth_wire[2] ),
	.cfg_devicewidth_wire_0(\c0|cfg_devicewidth_wire[0] ),
	.cfg_devicewidth_wire_1(\c0|cfg_devicewidth_wire[1] ),
	.cfg_devicewidth_wire_2(\c0|cfg_devicewidth_wire[2] ),
	.cfg_devicewidth_wire_3(\c0|cfg_devicewidth_wire[3] ),
	.cfg_interfacewidth_wire_0(\c0|cfg_interfacewidth_wire[0] ),
	.cfg_interfacewidth_wire_1(\c0|cfg_interfacewidth_wire[1] ),
	.cfg_interfacewidth_wire_2(\c0|cfg_interfacewidth_wire[2] ),
	.cfg_interfacewidth_wire_3(\c0|cfg_interfacewidth_wire[3] ),
	.cfg_interfacewidth_wire_4(\c0|cfg_interfacewidth_wire[4] ),
	.cfg_interfacewidth_wire_5(\c0|cfg_interfacewidth_wire[5] ),
	.cfg_interfacewidth_wire_6(\c0|cfg_interfacewidth_wire[6] ),
	.cfg_interfacewidth_wire_7(\c0|cfg_interfacewidth_wire[7] ),
	.cfg_rowaddrwidth_wire_0(\c0|cfg_rowaddrwidth_wire[0] ),
	.cfg_rowaddrwidth_wire_1(\c0|cfg_rowaddrwidth_wire[1] ),
	.cfg_rowaddrwidth_wire_2(\c0|cfg_rowaddrwidth_wire[2] ),
	.cfg_rowaddrwidth_wire_3(\c0|cfg_rowaddrwidth_wire[3] ),
	.cfg_rowaddrwidth_wire_4(\c0|cfg_rowaddrwidth_wire[4] ),
	.cfg_tcl_wire_0(\c0|cfg_tcl_wire[0] ),
	.cfg_tcl_wire_1(\c0|cfg_tcl_wire[1] ),
	.cfg_tcl_wire_2(\c0|cfg_tcl_wire[2] ),
	.cfg_tcl_wire_3(\c0|cfg_tcl_wire[3] ),
	.cfg_tcl_wire_4(\c0|cfg_tcl_wire[4] ),
	.cfg_tmrd_wire_0(\c0|cfg_tmrd_wire[0] ),
	.cfg_tmrd_wire_1(\c0|cfg_tmrd_wire[1] ),
	.cfg_tmrd_wire_2(\c0|cfg_tmrd_wire[2] ),
	.cfg_tmrd_wire_3(\c0|cfg_tmrd_wire[3] ),
	.cfg_trefi_wire_0(\c0|cfg_trefi_wire[0] ),
	.cfg_trefi_wire_1(\c0|cfg_trefi_wire[1] ),
	.cfg_trefi_wire_2(\c0|cfg_trefi_wire[2] ),
	.cfg_trefi_wire_3(\c0|cfg_trefi_wire[3] ),
	.cfg_trefi_wire_4(\c0|cfg_trefi_wire[4] ),
	.cfg_trefi_wire_5(\c0|cfg_trefi_wire[5] ),
	.cfg_trefi_wire_6(\c0|cfg_trefi_wire[6] ),
	.cfg_trefi_wire_7(\c0|cfg_trefi_wire[7] ),
	.cfg_trefi_wire_8(\c0|cfg_trefi_wire[8] ),
	.cfg_trefi_wire_9(\c0|cfg_trefi_wire[9] ),
	.cfg_trefi_wire_10(\c0|cfg_trefi_wire[10] ),
	.cfg_trefi_wire_11(\c0|cfg_trefi_wire[11] ),
	.cfg_trefi_wire_12(\c0|cfg_trefi_wire[12] ),
	.cfg_trfc_wire_0(\c0|cfg_trfc_wire[0] ),
	.cfg_trfc_wire_1(\c0|cfg_trfc_wire[1] ),
	.cfg_trfc_wire_2(\c0|cfg_trfc_wire[2] ),
	.cfg_trfc_wire_3(\c0|cfg_trfc_wire[3] ),
	.cfg_trfc_wire_4(\c0|cfg_trfc_wire[4] ),
	.cfg_trfc_wire_5(\c0|cfg_trfc_wire[5] ),
	.cfg_trfc_wire_6(\c0|cfg_trfc_wire[6] ),
	.cfg_trfc_wire_7(\c0|cfg_trfc_wire[7] ),
	.cfg_twr_wire_0(\c0|cfg_twr_wire[0] ),
	.cfg_twr_wire_1(\c0|cfg_twr_wire[1] ),
	.cfg_twr_wire_2(\c0|cfg_twr_wire[2] ),
	.cfg_twr_wire_3(\c0|cfg_twr_wire[3] ),
	.afi_mem_clk_disable_0(\c0|afi_mem_clk_disable[0] ),
	.cfg_dramconfig_wire_0(\c0|cfg_dramconfig_wire[0] ),
	.cfg_dramconfig_wire_1(\c0|cfg_dramconfig_wire[1] ),
	.cfg_dramconfig_wire_2(\c0|cfg_dramconfig_wire[2] ),
	.cfg_dramconfig_wire_3(\c0|cfg_dramconfig_wire[3] ),
	.cfg_dramconfig_wire_4(\c0|cfg_dramconfig_wire[4] ),
	.cfg_dramconfig_wire_5(\c0|cfg_dramconfig_wire[5] ),
	.cfg_dramconfig_wire_6(\c0|cfg_dramconfig_wire[6] ),
	.cfg_dramconfig_wire_7(\c0|cfg_dramconfig_wire[7] ),
	.cfg_dramconfig_wire_8(\c0|cfg_dramconfig_wire[8] ),
	.cfg_dramconfig_wire_9(\c0|cfg_dramconfig_wire[9] ),
	.cfg_dramconfig_wire_10(\c0|cfg_dramconfig_wire[10] ),
	.cfg_dramconfig_wire_11(\c0|cfg_dramconfig_wire[11] ),
	.cfg_dramconfig_wire_12(\c0|cfg_dramconfig_wire[12] ),
	.cfg_dramconfig_wire_13(\c0|cfg_dramconfig_wire[13] ),
	.cfg_dramconfig_wire_14(\c0|cfg_dramconfig_wire[14] ),
	.cfg_dramconfig_wire_15(\c0|cfg_dramconfig_wire[15] ),
	.cfg_dramconfig_wire_16(\c0|cfg_dramconfig_wire[16] ),
	.cfg_dramconfig_wire_17(\c0|cfg_dramconfig_wire[17] ),
	.cfg_dramconfig_wire_18(\c0|cfg_dramconfig_wire[18] ),
	.cfg_dramconfig_wire_19(\c0|cfg_dramconfig_wire[19] ),
	.cfg_dramconfig_wire_20(\c0|cfg_dramconfig_wire[20] ),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ),
	.dll_delayctrl_0(\dll|dll_delayctrl[0] ),
	.dll_delayctrl_1(\dll|dll_delayctrl[1] ),
	.dll_delayctrl_2(\dll|dll_delayctrl[2] ),
	.dll_delayctrl_3(\dll|dll_delayctrl[3] ),
	.dll_delayctrl_4(\dll|dll_delayctrl[4] ),
	.dll_delayctrl_5(\dll|dll_delayctrl[5] ),
	.dll_delayctrl_6(\dll|dll_delayctrl[6] ),
	.GND_port(GND_port));

Computer_System_hps_sdram_pll pll(
	.pll_mem_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ));

Computer_System_altera_mem_if_dll_cyclonev dll(
	.clk(\pll|pll_write_clk ),
	.dll_delayctrl({\dll|dll_delayctrl[6] ,\dll|dll_delayctrl[5] ,\dll|dll_delayctrl[4] ,\dll|dll_delayctrl[3] ,\dll|dll_delayctrl[2] ,\dll|dll_delayctrl[1] ,\dll|dll_delayctrl[0] }));

Computer_System_altera_mem_if_oct_cyclonev oct(
	.parallelterminationcontrol({parallelterminationcontrol_15,parallelterminationcontrol_14,parallelterminationcontrol_13,parallelterminationcontrol_12,parallelterminationcontrol_11,parallelterminationcontrol_10,parallelterminationcontrol_9,parallelterminationcontrol_8,
parallelterminationcontrol_7,parallelterminationcontrol_6,parallelterminationcontrol_5,parallelterminationcontrol_4,parallelterminationcontrol_3,parallelterminationcontrol_2,parallelterminationcontrol_1,parallelterminationcontrol_0}),
	.seriesterminationcontrol({seriesterminationcontrol_15,seriesterminationcontrol_14,seriesterminationcontrol_13,seriesterminationcontrol_12,seriesterminationcontrol_11,seriesterminationcontrol_10,seriesterminationcontrol_9,seriesterminationcontrol_8,seriesterminationcontrol_7,
seriesterminationcontrol_6,seriesterminationcontrol_5,seriesterminationcontrol_4,seriesterminationcontrol_3,seriesterminationcontrol_2,seriesterminationcontrol_1,seriesterminationcontrol_0}),
	.oct_rzqin(memory_oct_rzqin));

Computer_System_altera_mem_if_hard_memory_controller_top_cyclonev c0(
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid({\p0|umemphy|afi_rdata_valid[0] }),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata({\p0|umemphy|afi_rdata[79] ,\p0|umemphy|afi_rdata[78] ,\p0|umemphy|afi_rdata[77] ,\p0|umemphy|afi_rdata[76] ,\p0|umemphy|afi_rdata[75] ,\p0|umemphy|afi_rdata[74] ,\p0|umemphy|afi_rdata[73] ,\p0|umemphy|afi_rdata[72] ,\p0|umemphy|afi_rdata[71] ,
\p0|umemphy|afi_rdata[70] ,\p0|umemphy|afi_rdata[69] ,\p0|umemphy|afi_rdata[68] ,\p0|umemphy|afi_rdata[67] ,\p0|umemphy|afi_rdata[66] ,\p0|umemphy|afi_rdata[65] ,\p0|umemphy|afi_rdata[64] ,\p0|umemphy|afi_rdata[63] ,\p0|umemphy|afi_rdata[62] ,
\p0|umemphy|afi_rdata[61] ,\p0|umemphy|afi_rdata[60] ,\p0|umemphy|afi_rdata[59] ,\p0|umemphy|afi_rdata[58] ,\p0|umemphy|afi_rdata[57] ,\p0|umemphy|afi_rdata[56] ,\p0|umemphy|afi_rdata[55] ,\p0|umemphy|afi_rdata[54] ,\p0|umemphy|afi_rdata[53] ,
\p0|umemphy|afi_rdata[52] ,\p0|umemphy|afi_rdata[51] ,\p0|umemphy|afi_rdata[50] ,\p0|umemphy|afi_rdata[49] ,\p0|umemphy|afi_rdata[48] ,\p0|umemphy|afi_rdata[47] ,\p0|umemphy|afi_rdata[46] ,\p0|umemphy|afi_rdata[45] ,\p0|umemphy|afi_rdata[44] ,
\p0|umemphy|afi_rdata[43] ,\p0|umemphy|afi_rdata[42] ,\p0|umemphy|afi_rdata[41] ,\p0|umemphy|afi_rdata[40] ,\p0|umemphy|afi_rdata[39] ,\p0|umemphy|afi_rdata[38] ,\p0|umemphy|afi_rdata[37] ,\p0|umemphy|afi_rdata[36] ,\p0|umemphy|afi_rdata[35] ,
\p0|umemphy|afi_rdata[34] ,\p0|umemphy|afi_rdata[33] ,\p0|umemphy|afi_rdata[32] ,\p0|umemphy|afi_rdata[31] ,\p0|umemphy|afi_rdata[30] ,\p0|umemphy|afi_rdata[29] ,\p0|umemphy|afi_rdata[28] ,\p0|umemphy|afi_rdata[27] ,\p0|umemphy|afi_rdata[26] ,
\p0|umemphy|afi_rdata[25] ,\p0|umemphy|afi_rdata[24] ,\p0|umemphy|afi_rdata[23] ,\p0|umemphy|afi_rdata[22] ,\p0|umemphy|afi_rdata[21] ,\p0|umemphy|afi_rdata[20] ,\p0|umemphy|afi_rdata[19] ,\p0|umemphy|afi_rdata[18] ,\p0|umemphy|afi_rdata[17] ,
\p0|umemphy|afi_rdata[16] ,\p0|umemphy|afi_rdata[15] ,\p0|umemphy|afi_rdata[14] ,\p0|umemphy|afi_rdata[13] ,\p0|umemphy|afi_rdata[12] ,\p0|umemphy|afi_rdata[11] ,\p0|umemphy|afi_rdata[10] ,\p0|umemphy|afi_rdata[9] ,\p0|umemphy|afi_rdata[8] ,
\p0|umemphy|afi_rdata[7] ,\p0|umemphy|afi_rdata[6] ,\p0|umemphy|afi_rdata[5] ,\p0|umemphy|afi_rdata[4] ,\p0|umemphy|afi_rdata[3] ,\p0|umemphy|afi_rdata[2] ,\p0|umemphy|afi_rdata[1] ,\p0|umemphy|afi_rdata[0] }),
	.afi_wlat({\p0|umemphy|afi_wlat[3] ,\p0|umemphy|afi_wlat[2] ,\p0|umemphy|afi_wlat[1] ,\p0|umemphy|afi_wlat[0] }),
	.afi_cas_n({\c0|afi_cas_n[0] }),
	.afi_ras_n({\c0|afi_ras_n[0] }),
	.afi_rst_n({\c0|afi_rst_n[0] }),
	.afi_we_n({\c0|afi_we_n[0] }),
	.afi_addr({\c0|afi_addr[19] ,\c0|afi_addr[18] ,\c0|afi_addr[17] ,\c0|afi_addr[16] ,\c0|afi_addr[15] ,\c0|afi_addr[14] ,\c0|afi_addr[13] ,\c0|afi_addr[12] ,\c0|afi_addr[11] ,\c0|afi_addr[10] ,\c0|afi_addr[9] ,\c0|afi_addr[8] ,\c0|afi_addr[7] ,\c0|afi_addr[6] ,\c0|afi_addr[5] ,
\c0|afi_addr[4] ,\c0|afi_addr[3] ,\c0|afi_addr[2] ,\c0|afi_addr[1] ,\c0|afi_addr[0] }),
	.afi_ba({\c0|afi_ba[2] ,\c0|afi_ba[1] ,\c0|afi_ba[0] }),
	.afi_cke({\c0|afi_cke[1] ,\c0|afi_cke[0] }),
	.afi_cs_n({\c0|afi_cs_n[1] ,\c0|afi_cs_n[0] }),
	.afi_dm({\c0|afi_dm_int[9] ,\c0|afi_dm_int[8] ,\c0|afi_dm_int[7] ,\c0|afi_dm_int[6] ,\c0|afi_dm_int[5] ,\c0|afi_dm_int[4] ,\c0|afi_dm_int[3] ,\c0|afi_dm_int[2] ,\c0|afi_dm_int[1] ,\c0|afi_dm_int[0] }),
	.afi_dqs_burst({\c0|afi_dqs_burst[4] ,\c0|afi_dqs_burst[3] ,\c0|afi_dqs_burst[2] ,\c0|afi_dqs_burst[1] ,\c0|afi_dqs_burst[0] }),
	.afi_odt({\c0|afi_odt[1] ,\c0|afi_odt[0] }),
	.afi_rdata_en({\c0|afi_rdata_en[4] ,\c0|afi_rdata_en[3] ,\c0|afi_rdata_en[2] ,\c0|afi_rdata_en[1] ,\c0|afi_rdata_en[0] }),
	.afi_rdata_en_full({\c0|afi_rdata_en_full[4] ,\c0|afi_rdata_en_full[3] ,\c0|afi_rdata_en_full[2] ,\c0|afi_rdata_en_full[1] ,\c0|afi_rdata_en_full[0] }),
	.afi_wdata({\c0|afi_wdata_int[79] ,\c0|afi_wdata_int[78] ,\c0|afi_wdata_int[77] ,\c0|afi_wdata_int[76] ,\c0|afi_wdata_int[75] ,\c0|afi_wdata_int[74] ,\c0|afi_wdata_int[73] ,\c0|afi_wdata_int[72] ,\c0|afi_wdata_int[71] ,\c0|afi_wdata_int[70] ,\c0|afi_wdata_int[69] ,
\c0|afi_wdata_int[68] ,\c0|afi_wdata_int[67] ,\c0|afi_wdata_int[66] ,\c0|afi_wdata_int[65] ,\c0|afi_wdata_int[64] ,\c0|afi_wdata_int[63] ,\c0|afi_wdata_int[62] ,\c0|afi_wdata_int[61] ,\c0|afi_wdata_int[60] ,\c0|afi_wdata_int[59] ,\c0|afi_wdata_int[58] ,
\c0|afi_wdata_int[57] ,\c0|afi_wdata_int[56] ,\c0|afi_wdata_int[55] ,\c0|afi_wdata_int[54] ,\c0|afi_wdata_int[53] ,\c0|afi_wdata_int[52] ,\c0|afi_wdata_int[51] ,\c0|afi_wdata_int[50] ,\c0|afi_wdata_int[49] ,\c0|afi_wdata_int[48] ,\c0|afi_wdata_int[47] ,
\c0|afi_wdata_int[46] ,\c0|afi_wdata_int[45] ,\c0|afi_wdata_int[44] ,\c0|afi_wdata_int[43] ,\c0|afi_wdata_int[42] ,\c0|afi_wdata_int[41] ,\c0|afi_wdata_int[40] ,\c0|afi_wdata_int[39] ,\c0|afi_wdata_int[38] ,\c0|afi_wdata_int[37] ,\c0|afi_wdata_int[36] ,
\c0|afi_wdata_int[35] ,\c0|afi_wdata_int[34] ,\c0|afi_wdata_int[33] ,\c0|afi_wdata_int[32] ,\c0|afi_wdata_int[31] ,\c0|afi_wdata_int[30] ,\c0|afi_wdata_int[29] ,\c0|afi_wdata_int[28] ,\c0|afi_wdata_int[27] ,\c0|afi_wdata_int[26] ,\c0|afi_wdata_int[25] ,
\c0|afi_wdata_int[24] ,\c0|afi_wdata_int[23] ,\c0|afi_wdata_int[22] ,\c0|afi_wdata_int[21] ,\c0|afi_wdata_int[20] ,\c0|afi_wdata_int[19] ,\c0|afi_wdata_int[18] ,\c0|afi_wdata_int[17] ,\c0|afi_wdata_int[16] ,\c0|afi_wdata_int[15] ,\c0|afi_wdata_int[14] ,
\c0|afi_wdata_int[13] ,\c0|afi_wdata_int[12] ,\c0|afi_wdata_int[11] ,\c0|afi_wdata_int[10] ,\c0|afi_wdata_int[9] ,\c0|afi_wdata_int[8] ,\c0|afi_wdata_int[7] ,\c0|afi_wdata_int[6] ,\c0|afi_wdata_int[5] ,\c0|afi_wdata_int[4] ,\c0|afi_wdata_int[3] ,\c0|afi_wdata_int[2] ,
\c0|afi_wdata_int[1] ,\c0|afi_wdata_int[0] }),
	.afi_wdata_valid({\c0|afi_wdata_valid[4] ,\c0|afi_wdata_valid[3] ,\c0|afi_wdata_valid[2] ,\c0|afi_wdata_valid[1] ,\c0|afi_wdata_valid[0] }),
	.cfg_addlat({cfg_addlat_unconnected_wire_7,cfg_addlat_unconnected_wire_6,cfg_addlat_unconnected_wire_5,\c0|cfg_addlat_wire[4] ,\c0|cfg_addlat_wire[3] ,\c0|cfg_addlat_wire[2] ,\c0|cfg_addlat_wire[1] ,\c0|cfg_addlat_wire[0] }),
	.cfg_bankaddrwidth({cfg_bankaddrwidth_unconnected_wire_7,cfg_bankaddrwidth_unconnected_wire_6,cfg_bankaddrwidth_unconnected_wire_5,cfg_bankaddrwidth_unconnected_wire_4,cfg_bankaddrwidth_unconnected_wire_3,\c0|cfg_bankaddrwidth_wire[2] ,\c0|cfg_bankaddrwidth_wire[1] ,
\c0|cfg_bankaddrwidth_wire[0] }),
	.cfg_caswrlat({cfg_caswrlat_unconnected_wire_7,cfg_caswrlat_unconnected_wire_6,cfg_caswrlat_unconnected_wire_5,cfg_caswrlat_unconnected_wire_4,\c0|cfg_caswrlat_wire[3] ,\c0|cfg_caswrlat_wire[2] ,\c0|cfg_caswrlat_wire[1] ,\c0|cfg_caswrlat_wire[0] }),
	.cfg_coladdrwidth({cfg_coladdrwidth_unconnected_wire_7,cfg_coladdrwidth_unconnected_wire_6,cfg_coladdrwidth_unconnected_wire_5,\c0|cfg_coladdrwidth_wire[4] ,\c0|cfg_coladdrwidth_wire[3] ,\c0|cfg_coladdrwidth_wire[2] ,\c0|cfg_coladdrwidth_wire[1] ,\c0|cfg_coladdrwidth_wire[0] }),
	.cfg_csaddrwidth({cfg_csaddrwidth_unconnected_wire_7,cfg_csaddrwidth_unconnected_wire_6,cfg_csaddrwidth_unconnected_wire_5,cfg_csaddrwidth_unconnected_wire_4,cfg_csaddrwidth_unconnected_wire_3,\c0|cfg_csaddrwidth_wire[2] ,\c0|cfg_csaddrwidth_wire[1] ,\c0|cfg_csaddrwidth_wire[0] }),
	.cfg_devicewidth({cfg_devicewidth_unconnected_wire_7,cfg_devicewidth_unconnected_wire_6,cfg_devicewidth_unconnected_wire_5,cfg_devicewidth_unconnected_wire_4,\c0|cfg_devicewidth_wire[3] ,\c0|cfg_devicewidth_wire[2] ,\c0|cfg_devicewidth_wire[1] ,\c0|cfg_devicewidth_wire[0] }),
	.cfg_interfacewidth({\c0|cfg_interfacewidth_wire[7] ,\c0|cfg_interfacewidth_wire[6] ,\c0|cfg_interfacewidth_wire[5] ,\c0|cfg_interfacewidth_wire[4] ,\c0|cfg_interfacewidth_wire[3] ,\c0|cfg_interfacewidth_wire[2] ,\c0|cfg_interfacewidth_wire[1] ,\c0|cfg_interfacewidth_wire[0] }),
	.cfg_rowaddrwidth({cfg_rowaddrwidth_unconnected_wire_7,cfg_rowaddrwidth_unconnected_wire_6,cfg_rowaddrwidth_unconnected_wire_5,\c0|cfg_rowaddrwidth_wire[4] ,\c0|cfg_rowaddrwidth_wire[3] ,\c0|cfg_rowaddrwidth_wire[2] ,\c0|cfg_rowaddrwidth_wire[1] ,\c0|cfg_rowaddrwidth_wire[0] }),
	.cfg_tcl({cfg_tcl_unconnected_wire_7,cfg_tcl_unconnected_wire_6,cfg_tcl_unconnected_wire_5,\c0|cfg_tcl_wire[4] ,\c0|cfg_tcl_wire[3] ,\c0|cfg_tcl_wire[2] ,\c0|cfg_tcl_wire[1] ,\c0|cfg_tcl_wire[0] }),
	.cfg_tmrd({cfg_tmrd_unconnected_wire_7,cfg_tmrd_unconnected_wire_6,cfg_tmrd_unconnected_wire_5,cfg_tmrd_unconnected_wire_4,\c0|cfg_tmrd_wire[3] ,\c0|cfg_tmrd_wire[2] ,\c0|cfg_tmrd_wire[1] ,\c0|cfg_tmrd_wire[0] }),
	.cfg_trefi({cfg_trefi_unconnected_wire_15,cfg_trefi_unconnected_wire_14,cfg_trefi_unconnected_wire_13,\c0|cfg_trefi_wire[12] ,\c0|cfg_trefi_wire[11] ,\c0|cfg_trefi_wire[10] ,\c0|cfg_trefi_wire[9] ,\c0|cfg_trefi_wire[8] ,\c0|cfg_trefi_wire[7] ,\c0|cfg_trefi_wire[6] ,
\c0|cfg_trefi_wire[5] ,\c0|cfg_trefi_wire[4] ,\c0|cfg_trefi_wire[3] ,\c0|cfg_trefi_wire[2] ,\c0|cfg_trefi_wire[1] ,\c0|cfg_trefi_wire[0] }),
	.cfg_trfc({\c0|cfg_trfc_wire[7] ,\c0|cfg_trfc_wire[6] ,\c0|cfg_trfc_wire[5] ,\c0|cfg_trfc_wire[4] ,\c0|cfg_trfc_wire[3] ,\c0|cfg_trfc_wire[2] ,\c0|cfg_trfc_wire[1] ,\c0|cfg_trfc_wire[0] }),
	.cfg_twr({cfg_twr_unconnected_wire_7,cfg_twr_unconnected_wire_6,cfg_twr_unconnected_wire_5,cfg_twr_unconnected_wire_4,\c0|cfg_twr_wire[3] ,\c0|cfg_twr_wire[2] ,\c0|cfg_twr_wire[1] ,\c0|cfg_twr_wire[0] }),
	.afi_mem_clk_disable({\c0|afi_mem_clk_disable[0] }),
	.cfg_dramconfig({cfg_dramconfig_unconnected_wire_23,cfg_dramconfig_unconnected_wire_22,cfg_dramconfig_unconnected_wire_21,\c0|cfg_dramconfig_wire[20] ,\c0|cfg_dramconfig_wire[19] ,\c0|cfg_dramconfig_wire[18] ,\c0|cfg_dramconfig_wire[17] ,\c0|cfg_dramconfig_wire[16] ,
\c0|cfg_dramconfig_wire[15] ,\c0|cfg_dramconfig_wire[14] ,\c0|cfg_dramconfig_wire[13] ,\c0|cfg_dramconfig_wire[12] ,\c0|cfg_dramconfig_wire[11] ,\c0|cfg_dramconfig_wire[10] ,\c0|cfg_dramconfig_wire[9] ,\c0|cfg_dramconfig_wire[8] ,\c0|cfg_dramconfig_wire[7] ,
\c0|cfg_dramconfig_wire[6] ,\c0|cfg_dramconfig_wire[5] ,\c0|cfg_dramconfig_wire[4] ,\c0|cfg_dramconfig_wire[3] ,\c0|cfg_dramconfig_wire[2] ,\c0|cfg_dramconfig_wire[1] ,\c0|cfg_dramconfig_wire[0] }),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ));

endmodule

module Computer_System_altera_mem_if_dll_cyclonev (
	clk,
	dll_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	[6:0] dll_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [6:0] dll_wys_m_DELAYCTRLOUT_bus;

assign dll_delayctrl[0] = dll_wys_m_DELAYCTRLOUT_bus[0];
assign dll_delayctrl[1] = dll_wys_m_DELAYCTRLOUT_bus[1];
assign dll_delayctrl[2] = dll_wys_m_DELAYCTRLOUT_bus[2];
assign dll_delayctrl[3] = dll_wys_m_DELAYCTRLOUT_bus[3];
assign dll_delayctrl[4] = dll_wys_m_DELAYCTRLOUT_bus[4];
assign dll_delayctrl[5] = dll_wys_m_DELAYCTRLOUT_bus[5];
assign dll_delayctrl[6] = dll_wys_m_DELAYCTRLOUT_bus[6];

cyclonev_dll dll_wys_m(
	.clk(clk),
	.aload(vcc),
	.upndnin(gnd),
	.upndninclkena(gnd),
	.dqsupdate(),
	.upndnout(),
	.delayctrlout(dll_wys_m_DELAYCTRLOUT_bus));
defparam dll_wys_m.delayctrlout_mode = "normal";
defparam dll_wys_m.input_frequency = "2500 ps";
defparam dll_wys_m.jitter_reduction = "true";
defparam dll_wys_m.sim_buffer_delay_increment = 10;
defparam dll_wys_m.sim_buffer_intrinsic_delay = 175;
defparam dll_wys_m.sim_valid_lock = 16;
defparam dll_wys_m.sim_valid_lockcount = 0;
defparam dll_wys_m.static_delay_ctrl = 8;
defparam dll_wys_m.upndnout_mode = "clock";
defparam dll_wys_m.use_upndnin = "false";
defparam dll_wys_m.use_upndninclkena = "false";

endmodule

module Computer_System_altera_mem_if_hard_memory_controller_top_cyclonev (
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk)/* synthesis synthesis_greybox=0 */;
input 	afi_cal_fail;
input 	afi_cal_success;
input 	[0:0] afi_rdata_valid;
input 	ctl_reset_n;
input 	[79:0] afi_rdata;
input 	[3:0] afi_wlat;
output 	[0:0] afi_cas_n;
output 	[0:0] afi_ras_n;
output 	[0:0] afi_rst_n;
output 	[0:0] afi_we_n;
output 	[19:0] afi_addr;
output 	[2:0] afi_ba;
output 	[1:0] afi_cke;
output 	[1:0] afi_cs_n;
output 	[9:0] afi_dm;
output 	[4:0] afi_dqs_burst;
output 	[1:0] afi_odt;
output 	[4:0] afi_rdata_en;
output 	[4:0] afi_rdata_en_full;
output 	[79:0] afi_wdata;
output 	[4:0] afi_wdata_valid;
output 	[7:0] cfg_addlat;
output 	[7:0] cfg_bankaddrwidth;
output 	[7:0] cfg_caswrlat;
output 	[7:0] cfg_coladdrwidth;
output 	[7:0] cfg_csaddrwidth;
output 	[7:0] cfg_devicewidth;
output 	[7:0] cfg_interfacewidth;
output 	[7:0] cfg_rowaddrwidth;
output 	[7:0] cfg_tcl;
output 	[7:0] cfg_tmrd;
output 	[15:0] cfg_trefi;
output 	[7:0] cfg_trfc;
output 	[7:0] cfg_twr;
output 	[0:0] afi_mem_clk_disable;
output 	[23:0] cfg_dramconfig;
input 	ctl_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [19:0] hmc_inst_AFIADDR_bus;
wire [2:0] hmc_inst_AFIBA_bus;
wire [1:0] hmc_inst_AFICKE_bus;
wire [1:0] hmc_inst_AFICSN_bus;
wire [9:0] hmc_inst_AFIDM_bus;
wire [4:0] hmc_inst_AFIDQSBURST_bus;
wire [1:0] hmc_inst_AFIODT_bus;
wire [4:0] hmc_inst_AFIRDATAEN_bus;
wire [4:0] hmc_inst_AFIRDATAENFULL_bus;
wire [79:0] hmc_inst_AFIWDATA_bus;
wire [4:0] hmc_inst_AFIWDATAVALID_bus;
wire [4:0] hmc_inst_CFGADDLAT_bus;
wire [2:0] hmc_inst_CFGBANKADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGCASWRLAT_bus;
wire [4:0] hmc_inst_CFGCOLADDRWIDTH_bus;
wire [2:0] hmc_inst_CFGCSADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGDEVICEWIDTH_bus;
wire [7:0] hmc_inst_CFGINTERFACEWIDTH_bus;
wire [4:0] hmc_inst_CFGROWADDRWIDTH_bus;
wire [4:0] hmc_inst_CFGTCL_bus;
wire [3:0] hmc_inst_CFGTMRD_bus;
wire [12:0] hmc_inst_CFGTREFI_bus;
wire [7:0] hmc_inst_CFGTRFC_bus;
wire [3:0] hmc_inst_CFGTWR_bus;
wire [1:0] hmc_inst_CTLMEMCLKDISABLE_bus;
wire [20:0] hmc_inst_DRAMCONFIG_bus;

assign afi_addr[0] = hmc_inst_AFIADDR_bus[0];
assign afi_addr[1] = hmc_inst_AFIADDR_bus[1];
assign afi_addr[2] = hmc_inst_AFIADDR_bus[2];
assign afi_addr[3] = hmc_inst_AFIADDR_bus[3];
assign afi_addr[4] = hmc_inst_AFIADDR_bus[4];
assign afi_addr[5] = hmc_inst_AFIADDR_bus[5];
assign afi_addr[6] = hmc_inst_AFIADDR_bus[6];
assign afi_addr[7] = hmc_inst_AFIADDR_bus[7];
assign afi_addr[8] = hmc_inst_AFIADDR_bus[8];
assign afi_addr[9] = hmc_inst_AFIADDR_bus[9];
assign afi_addr[10] = hmc_inst_AFIADDR_bus[10];
assign afi_addr[11] = hmc_inst_AFIADDR_bus[11];
assign afi_addr[12] = hmc_inst_AFIADDR_bus[12];
assign afi_addr[13] = hmc_inst_AFIADDR_bus[13];
assign afi_addr[14] = hmc_inst_AFIADDR_bus[14];
assign afi_addr[15] = hmc_inst_AFIADDR_bus[15];
assign afi_addr[16] = hmc_inst_AFIADDR_bus[16];
assign afi_addr[17] = hmc_inst_AFIADDR_bus[17];
assign afi_addr[18] = hmc_inst_AFIADDR_bus[18];
assign afi_addr[19] = hmc_inst_AFIADDR_bus[19];

assign afi_ba[0] = hmc_inst_AFIBA_bus[0];
assign afi_ba[1] = hmc_inst_AFIBA_bus[1];
assign afi_ba[2] = hmc_inst_AFIBA_bus[2];

assign afi_cke[0] = hmc_inst_AFICKE_bus[0];
assign afi_cke[1] = hmc_inst_AFICKE_bus[1];

assign afi_cs_n[0] = hmc_inst_AFICSN_bus[0];
assign afi_cs_n[1] = hmc_inst_AFICSN_bus[1];

assign afi_dm[0] = hmc_inst_AFIDM_bus[0];
assign afi_dm[1] = hmc_inst_AFIDM_bus[1];
assign afi_dm[2] = hmc_inst_AFIDM_bus[2];
assign afi_dm[3] = hmc_inst_AFIDM_bus[3];
assign afi_dm[4] = hmc_inst_AFIDM_bus[4];
assign afi_dm[5] = hmc_inst_AFIDM_bus[5];
assign afi_dm[6] = hmc_inst_AFIDM_bus[6];
assign afi_dm[7] = hmc_inst_AFIDM_bus[7];
assign afi_dm[8] = hmc_inst_AFIDM_bus[8];
assign afi_dm[9] = hmc_inst_AFIDM_bus[9];

assign afi_dqs_burst[0] = hmc_inst_AFIDQSBURST_bus[0];
assign afi_dqs_burst[1] = hmc_inst_AFIDQSBURST_bus[1];
assign afi_dqs_burst[2] = hmc_inst_AFIDQSBURST_bus[2];
assign afi_dqs_burst[3] = hmc_inst_AFIDQSBURST_bus[3];
assign afi_dqs_burst[4] = hmc_inst_AFIDQSBURST_bus[4];

assign afi_odt[0] = hmc_inst_AFIODT_bus[0];
assign afi_odt[1] = hmc_inst_AFIODT_bus[1];

assign afi_rdata_en[0] = hmc_inst_AFIRDATAEN_bus[0];
assign afi_rdata_en[1] = hmc_inst_AFIRDATAEN_bus[1];
assign afi_rdata_en[2] = hmc_inst_AFIRDATAEN_bus[2];
assign afi_rdata_en[3] = hmc_inst_AFIRDATAEN_bus[3];
assign afi_rdata_en[4] = hmc_inst_AFIRDATAEN_bus[4];

assign afi_rdata_en_full[0] = hmc_inst_AFIRDATAENFULL_bus[0];
assign afi_rdata_en_full[1] = hmc_inst_AFIRDATAENFULL_bus[1];
assign afi_rdata_en_full[2] = hmc_inst_AFIRDATAENFULL_bus[2];
assign afi_rdata_en_full[3] = hmc_inst_AFIRDATAENFULL_bus[3];
assign afi_rdata_en_full[4] = hmc_inst_AFIRDATAENFULL_bus[4];

assign afi_wdata[0] = hmc_inst_AFIWDATA_bus[0];
assign afi_wdata[1] = hmc_inst_AFIWDATA_bus[1];
assign afi_wdata[2] = hmc_inst_AFIWDATA_bus[2];
assign afi_wdata[3] = hmc_inst_AFIWDATA_bus[3];
assign afi_wdata[4] = hmc_inst_AFIWDATA_bus[4];
assign afi_wdata[5] = hmc_inst_AFIWDATA_bus[5];
assign afi_wdata[6] = hmc_inst_AFIWDATA_bus[6];
assign afi_wdata[7] = hmc_inst_AFIWDATA_bus[7];
assign afi_wdata[8] = hmc_inst_AFIWDATA_bus[8];
assign afi_wdata[9] = hmc_inst_AFIWDATA_bus[9];
assign afi_wdata[10] = hmc_inst_AFIWDATA_bus[10];
assign afi_wdata[11] = hmc_inst_AFIWDATA_bus[11];
assign afi_wdata[12] = hmc_inst_AFIWDATA_bus[12];
assign afi_wdata[13] = hmc_inst_AFIWDATA_bus[13];
assign afi_wdata[14] = hmc_inst_AFIWDATA_bus[14];
assign afi_wdata[15] = hmc_inst_AFIWDATA_bus[15];
assign afi_wdata[16] = hmc_inst_AFIWDATA_bus[16];
assign afi_wdata[17] = hmc_inst_AFIWDATA_bus[17];
assign afi_wdata[18] = hmc_inst_AFIWDATA_bus[18];
assign afi_wdata[19] = hmc_inst_AFIWDATA_bus[19];
assign afi_wdata[20] = hmc_inst_AFIWDATA_bus[20];
assign afi_wdata[21] = hmc_inst_AFIWDATA_bus[21];
assign afi_wdata[22] = hmc_inst_AFIWDATA_bus[22];
assign afi_wdata[23] = hmc_inst_AFIWDATA_bus[23];
assign afi_wdata[24] = hmc_inst_AFIWDATA_bus[24];
assign afi_wdata[25] = hmc_inst_AFIWDATA_bus[25];
assign afi_wdata[26] = hmc_inst_AFIWDATA_bus[26];
assign afi_wdata[27] = hmc_inst_AFIWDATA_bus[27];
assign afi_wdata[28] = hmc_inst_AFIWDATA_bus[28];
assign afi_wdata[29] = hmc_inst_AFIWDATA_bus[29];
assign afi_wdata[30] = hmc_inst_AFIWDATA_bus[30];
assign afi_wdata[31] = hmc_inst_AFIWDATA_bus[31];
assign afi_wdata[32] = hmc_inst_AFIWDATA_bus[32];
assign afi_wdata[33] = hmc_inst_AFIWDATA_bus[33];
assign afi_wdata[34] = hmc_inst_AFIWDATA_bus[34];
assign afi_wdata[35] = hmc_inst_AFIWDATA_bus[35];
assign afi_wdata[36] = hmc_inst_AFIWDATA_bus[36];
assign afi_wdata[37] = hmc_inst_AFIWDATA_bus[37];
assign afi_wdata[38] = hmc_inst_AFIWDATA_bus[38];
assign afi_wdata[39] = hmc_inst_AFIWDATA_bus[39];
assign afi_wdata[40] = hmc_inst_AFIWDATA_bus[40];
assign afi_wdata[41] = hmc_inst_AFIWDATA_bus[41];
assign afi_wdata[42] = hmc_inst_AFIWDATA_bus[42];
assign afi_wdata[43] = hmc_inst_AFIWDATA_bus[43];
assign afi_wdata[44] = hmc_inst_AFIWDATA_bus[44];
assign afi_wdata[45] = hmc_inst_AFIWDATA_bus[45];
assign afi_wdata[46] = hmc_inst_AFIWDATA_bus[46];
assign afi_wdata[47] = hmc_inst_AFIWDATA_bus[47];
assign afi_wdata[48] = hmc_inst_AFIWDATA_bus[48];
assign afi_wdata[49] = hmc_inst_AFIWDATA_bus[49];
assign afi_wdata[50] = hmc_inst_AFIWDATA_bus[50];
assign afi_wdata[51] = hmc_inst_AFIWDATA_bus[51];
assign afi_wdata[52] = hmc_inst_AFIWDATA_bus[52];
assign afi_wdata[53] = hmc_inst_AFIWDATA_bus[53];
assign afi_wdata[54] = hmc_inst_AFIWDATA_bus[54];
assign afi_wdata[55] = hmc_inst_AFIWDATA_bus[55];
assign afi_wdata[56] = hmc_inst_AFIWDATA_bus[56];
assign afi_wdata[57] = hmc_inst_AFIWDATA_bus[57];
assign afi_wdata[58] = hmc_inst_AFIWDATA_bus[58];
assign afi_wdata[59] = hmc_inst_AFIWDATA_bus[59];
assign afi_wdata[60] = hmc_inst_AFIWDATA_bus[60];
assign afi_wdata[61] = hmc_inst_AFIWDATA_bus[61];
assign afi_wdata[62] = hmc_inst_AFIWDATA_bus[62];
assign afi_wdata[63] = hmc_inst_AFIWDATA_bus[63];
assign afi_wdata[64] = hmc_inst_AFIWDATA_bus[64];
assign afi_wdata[65] = hmc_inst_AFIWDATA_bus[65];
assign afi_wdata[66] = hmc_inst_AFIWDATA_bus[66];
assign afi_wdata[67] = hmc_inst_AFIWDATA_bus[67];
assign afi_wdata[68] = hmc_inst_AFIWDATA_bus[68];
assign afi_wdata[69] = hmc_inst_AFIWDATA_bus[69];
assign afi_wdata[70] = hmc_inst_AFIWDATA_bus[70];
assign afi_wdata[71] = hmc_inst_AFIWDATA_bus[71];
assign afi_wdata[72] = hmc_inst_AFIWDATA_bus[72];
assign afi_wdata[73] = hmc_inst_AFIWDATA_bus[73];
assign afi_wdata[74] = hmc_inst_AFIWDATA_bus[74];
assign afi_wdata[75] = hmc_inst_AFIWDATA_bus[75];
assign afi_wdata[76] = hmc_inst_AFIWDATA_bus[76];
assign afi_wdata[77] = hmc_inst_AFIWDATA_bus[77];
assign afi_wdata[78] = hmc_inst_AFIWDATA_bus[78];
assign afi_wdata[79] = hmc_inst_AFIWDATA_bus[79];

assign afi_wdata_valid[0] = hmc_inst_AFIWDATAVALID_bus[0];
assign afi_wdata_valid[1] = hmc_inst_AFIWDATAVALID_bus[1];
assign afi_wdata_valid[2] = hmc_inst_AFIWDATAVALID_bus[2];
assign afi_wdata_valid[3] = hmc_inst_AFIWDATAVALID_bus[3];
assign afi_wdata_valid[4] = hmc_inst_AFIWDATAVALID_bus[4];

assign cfg_addlat[0] = hmc_inst_CFGADDLAT_bus[0];
assign cfg_addlat[1] = hmc_inst_CFGADDLAT_bus[1];
assign cfg_addlat[2] = hmc_inst_CFGADDLAT_bus[2];
assign cfg_addlat[3] = hmc_inst_CFGADDLAT_bus[3];
assign cfg_addlat[4] = hmc_inst_CFGADDLAT_bus[4];

assign cfg_bankaddrwidth[0] = hmc_inst_CFGBANKADDRWIDTH_bus[0];
assign cfg_bankaddrwidth[1] = hmc_inst_CFGBANKADDRWIDTH_bus[1];
assign cfg_bankaddrwidth[2] = hmc_inst_CFGBANKADDRWIDTH_bus[2];

assign cfg_caswrlat[0] = hmc_inst_CFGCASWRLAT_bus[0];
assign cfg_caswrlat[1] = hmc_inst_CFGCASWRLAT_bus[1];
assign cfg_caswrlat[2] = hmc_inst_CFGCASWRLAT_bus[2];
assign cfg_caswrlat[3] = hmc_inst_CFGCASWRLAT_bus[3];

assign cfg_coladdrwidth[0] = hmc_inst_CFGCOLADDRWIDTH_bus[0];
assign cfg_coladdrwidth[1] = hmc_inst_CFGCOLADDRWIDTH_bus[1];
assign cfg_coladdrwidth[2] = hmc_inst_CFGCOLADDRWIDTH_bus[2];
assign cfg_coladdrwidth[3] = hmc_inst_CFGCOLADDRWIDTH_bus[3];
assign cfg_coladdrwidth[4] = hmc_inst_CFGCOLADDRWIDTH_bus[4];

assign cfg_csaddrwidth[0] = hmc_inst_CFGCSADDRWIDTH_bus[0];
assign cfg_csaddrwidth[1] = hmc_inst_CFGCSADDRWIDTH_bus[1];
assign cfg_csaddrwidth[2] = hmc_inst_CFGCSADDRWIDTH_bus[2];

assign cfg_devicewidth[0] = hmc_inst_CFGDEVICEWIDTH_bus[0];
assign cfg_devicewidth[1] = hmc_inst_CFGDEVICEWIDTH_bus[1];
assign cfg_devicewidth[2] = hmc_inst_CFGDEVICEWIDTH_bus[2];
assign cfg_devicewidth[3] = hmc_inst_CFGDEVICEWIDTH_bus[3];

assign cfg_interfacewidth[0] = hmc_inst_CFGINTERFACEWIDTH_bus[0];
assign cfg_interfacewidth[1] = hmc_inst_CFGINTERFACEWIDTH_bus[1];
assign cfg_interfacewidth[2] = hmc_inst_CFGINTERFACEWIDTH_bus[2];
assign cfg_interfacewidth[3] = hmc_inst_CFGINTERFACEWIDTH_bus[3];
assign cfg_interfacewidth[4] = hmc_inst_CFGINTERFACEWIDTH_bus[4];
assign cfg_interfacewidth[5] = hmc_inst_CFGINTERFACEWIDTH_bus[5];
assign cfg_interfacewidth[6] = hmc_inst_CFGINTERFACEWIDTH_bus[6];
assign cfg_interfacewidth[7] = hmc_inst_CFGINTERFACEWIDTH_bus[7];

assign cfg_rowaddrwidth[0] = hmc_inst_CFGROWADDRWIDTH_bus[0];
assign cfg_rowaddrwidth[1] = hmc_inst_CFGROWADDRWIDTH_bus[1];
assign cfg_rowaddrwidth[2] = hmc_inst_CFGROWADDRWIDTH_bus[2];
assign cfg_rowaddrwidth[3] = hmc_inst_CFGROWADDRWIDTH_bus[3];
assign cfg_rowaddrwidth[4] = hmc_inst_CFGROWADDRWIDTH_bus[4];

assign cfg_tcl[0] = hmc_inst_CFGTCL_bus[0];
assign cfg_tcl[1] = hmc_inst_CFGTCL_bus[1];
assign cfg_tcl[2] = hmc_inst_CFGTCL_bus[2];
assign cfg_tcl[3] = hmc_inst_CFGTCL_bus[3];
assign cfg_tcl[4] = hmc_inst_CFGTCL_bus[4];

assign cfg_tmrd[0] = hmc_inst_CFGTMRD_bus[0];
assign cfg_tmrd[1] = hmc_inst_CFGTMRD_bus[1];
assign cfg_tmrd[2] = hmc_inst_CFGTMRD_bus[2];
assign cfg_tmrd[3] = hmc_inst_CFGTMRD_bus[3];

assign cfg_trefi[0] = hmc_inst_CFGTREFI_bus[0];
assign cfg_trefi[1] = hmc_inst_CFGTREFI_bus[1];
assign cfg_trefi[2] = hmc_inst_CFGTREFI_bus[2];
assign cfg_trefi[3] = hmc_inst_CFGTREFI_bus[3];
assign cfg_trefi[4] = hmc_inst_CFGTREFI_bus[4];
assign cfg_trefi[5] = hmc_inst_CFGTREFI_bus[5];
assign cfg_trefi[6] = hmc_inst_CFGTREFI_bus[6];
assign cfg_trefi[7] = hmc_inst_CFGTREFI_bus[7];
assign cfg_trefi[8] = hmc_inst_CFGTREFI_bus[8];
assign cfg_trefi[9] = hmc_inst_CFGTREFI_bus[9];
assign cfg_trefi[10] = hmc_inst_CFGTREFI_bus[10];
assign cfg_trefi[11] = hmc_inst_CFGTREFI_bus[11];
assign cfg_trefi[12] = hmc_inst_CFGTREFI_bus[12];

assign cfg_trfc[0] = hmc_inst_CFGTRFC_bus[0];
assign cfg_trfc[1] = hmc_inst_CFGTRFC_bus[1];
assign cfg_trfc[2] = hmc_inst_CFGTRFC_bus[2];
assign cfg_trfc[3] = hmc_inst_CFGTRFC_bus[3];
assign cfg_trfc[4] = hmc_inst_CFGTRFC_bus[4];
assign cfg_trfc[5] = hmc_inst_CFGTRFC_bus[5];
assign cfg_trfc[6] = hmc_inst_CFGTRFC_bus[6];
assign cfg_trfc[7] = hmc_inst_CFGTRFC_bus[7];

assign cfg_twr[0] = hmc_inst_CFGTWR_bus[0];
assign cfg_twr[1] = hmc_inst_CFGTWR_bus[1];
assign cfg_twr[2] = hmc_inst_CFGTWR_bus[2];
assign cfg_twr[3] = hmc_inst_CFGTWR_bus[3];

assign afi_mem_clk_disable[0] = hmc_inst_CTLMEMCLKDISABLE_bus[0];

assign cfg_dramconfig[0] = hmc_inst_DRAMCONFIG_bus[0];
assign cfg_dramconfig[1] = hmc_inst_DRAMCONFIG_bus[1];
assign cfg_dramconfig[2] = hmc_inst_DRAMCONFIG_bus[2];
assign cfg_dramconfig[3] = hmc_inst_DRAMCONFIG_bus[3];
assign cfg_dramconfig[4] = hmc_inst_DRAMCONFIG_bus[4];
assign cfg_dramconfig[5] = hmc_inst_DRAMCONFIG_bus[5];
assign cfg_dramconfig[6] = hmc_inst_DRAMCONFIG_bus[6];
assign cfg_dramconfig[7] = hmc_inst_DRAMCONFIG_bus[7];
assign cfg_dramconfig[8] = hmc_inst_DRAMCONFIG_bus[8];
assign cfg_dramconfig[9] = hmc_inst_DRAMCONFIG_bus[9];
assign cfg_dramconfig[10] = hmc_inst_DRAMCONFIG_bus[10];
assign cfg_dramconfig[11] = hmc_inst_DRAMCONFIG_bus[11];
assign cfg_dramconfig[12] = hmc_inst_DRAMCONFIG_bus[12];
assign cfg_dramconfig[13] = hmc_inst_DRAMCONFIG_bus[13];
assign cfg_dramconfig[14] = hmc_inst_DRAMCONFIG_bus[14];
assign cfg_dramconfig[15] = hmc_inst_DRAMCONFIG_bus[15];
assign cfg_dramconfig[16] = hmc_inst_DRAMCONFIG_bus[16];
assign cfg_dramconfig[17] = hmc_inst_DRAMCONFIG_bus[17];
assign cfg_dramconfig[18] = hmc_inst_DRAMCONFIG_bus[18];
assign cfg_dramconfig[19] = hmc_inst_DRAMCONFIG_bus[19];
assign cfg_dramconfig[20] = hmc_inst_DRAMCONFIG_bus[20];

cyclonev_hmc hmc_inst(
	.afirdatavalid(afi_rdata_valid[0]),
	.csrclk(gnd),
	.csrdin(gnd),
	.csren(gnd),
	.ctlcalfail(afi_cal_fail),
	.ctlcalsuccess(afi_cal_success),
	.ctlclk(ctl_clk),
	.ctlresetn(ctl_reset_n),
	.globalresetn(gnd),
	.iavstcmdresetn0(vcc),
	.iavstcmdresetn1(vcc),
	.iavstcmdresetn2(vcc),
	.iavstcmdresetn3(vcc),
	.iavstcmdresetn4(vcc),
	.iavstcmdresetn5(vcc),
	.iavstrdclk0(gnd),
	.iavstrdclk1(gnd),
	.iavstrdclk2(gnd),
	.iavstrdclk3(gnd),
	.iavstrdready0(vcc),
	.iavstrdready1(vcc),
	.iavstrdready2(vcc),
	.iavstrdready3(vcc),
	.iavstrdresetn0(vcc),
	.iavstrdresetn1(vcc),
	.iavstrdresetn2(vcc),
	.iavstrdresetn3(vcc),
	.iavstwrackready0(vcc),
	.iavstwrackready1(vcc),
	.iavstwrackready2(vcc),
	.iavstwrackready3(vcc),
	.iavstwrackready4(vcc),
	.iavstwrackready5(vcc),
	.iavstwrclk0(gnd),
	.iavstwrclk1(gnd),
	.iavstwrclk2(gnd),
	.iavstwrclk3(gnd),
	.iavstwrresetn0(vcc),
	.iavstwrresetn1(vcc),
	.iavstwrresetn2(vcc),
	.iavstwrresetn3(vcc),
	.localdeeppowerdnreq(gnd),
	.localrefreshreq(gnd),
	.localselfrfshreq(gnd),
	.mmrbe(gnd),
	.mmrburstbegin(vcc),
	.mmrclk(gnd),
	.mmrreadreq(gnd),
	.mmrresetn(vcc),
	.mmrwritereq(gnd),
	.portclk0(gnd),
	.portclk1(gnd),
	.portclk2(gnd),
	.portclk3(gnd),
	.portclk4(gnd),
	.portclk5(gnd),
	.scanenable(gnd),
	.scbe(gnd),
	.scburstbegin(gnd),
	.scclk(gnd),
	.screadreq(gnd),
	.scresetn(vcc),
	.scwritereq(gnd),
	.afirdata({afi_rdata[79],afi_rdata[78],afi_rdata[77],afi_rdata[76],afi_rdata[75],afi_rdata[74],afi_rdata[73],afi_rdata[72],afi_rdata[71],afi_rdata[70],afi_rdata[69],afi_rdata[68],afi_rdata[67],afi_rdata[66],afi_rdata[65],afi_rdata[64],afi_rdata[63],afi_rdata[62],afi_rdata[61],afi_rdata[60],afi_rdata[59],afi_rdata[58],afi_rdata[57],afi_rdata[56],afi_rdata[55],afi_rdata[54],afi_rdata[53],afi_rdata[52],
afi_rdata[51],afi_rdata[50],afi_rdata[49],afi_rdata[48],afi_rdata[47],afi_rdata[46],afi_rdata[45],afi_rdata[44],afi_rdata[43],afi_rdata[42],afi_rdata[41],afi_rdata[40],afi_rdata[39],afi_rdata[38],afi_rdata[37],afi_rdata[36],afi_rdata[35],afi_rdata[34],afi_rdata[33],afi_rdata[32],afi_rdata[31],afi_rdata[30],afi_rdata[29],afi_rdata[28],afi_rdata[27],afi_rdata[26],afi_rdata[25],afi_rdata[24],
afi_rdata[23],afi_rdata[22],afi_rdata[21],afi_rdata[20],afi_rdata[19],afi_rdata[18],afi_rdata[17],afi_rdata[16],afi_rdata[15],afi_rdata[14],afi_rdata[13],afi_rdata[12],afi_rdata[11],afi_rdata[10],afi_rdata[9],afi_rdata[8],afi_rdata[7],afi_rdata[6],afi_rdata[5],afi_rdata[4],afi_rdata[3],afi_rdata[2],afi_rdata[1],afi_rdata[0]}),
	.afiseqbusy({gnd,gnd}),
	.afiwlat({afi_wlat[3],afi_wlat[2],afi_wlat[1],afi_wlat[0]}),
	.bondingin1({gnd,gnd,gnd,gnd}),
	.bondingin2({gnd,gnd,gnd,gnd,gnd,gnd}),
	.bondingin3({gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata4({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata5({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.localdeeppowerdnchip({gnd,gnd}),
	.localrefreshchip({gnd,gnd}),
	.localselfrfshchip({gnd,gnd}),
	.mmraddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.mmrburstcount({gnd,vcc}),
	.mmrwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scburstcount({gnd,gnd}),
	.scwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.aficasn(afi_cas_n[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.csrdout(),
	.ctlcalreq(),
	.ctlinitreq(),
	.localdeeppowerdnack(),
	.localinitdone(),
	.localpowerdownack(),
	.localrefreshack(),
	.localselfrfshack(),
	.localstsctlempty(),
	.mmrrdatavalid(),
	.mmrwaitrequest(),
	.oammready0(),
	.oammready1(),
	.oammready2(),
	.oammready3(),
	.oammready4(),
	.oammready5(),
	.ordavstvalid0(),
	.ordavstvalid1(),
	.ordavstvalid2(),
	.ordavstvalid3(),
	.owrackavstdata0(),
	.owrackavstdata1(),
	.owrackavstdata2(),
	.owrackavstdata3(),
	.owrackavstdata4(),
	.owrackavstdata5(),
	.owrackavstvalid0(),
	.owrackavstvalid1(),
	.owrackavstvalid2(),
	.owrackavstvalid3(),
	.owrackavstvalid4(),
	.owrackavstvalid5(),
	.scrdatavalid(),
	.scwaitrequest(),
	.afiaddr(hmc_inst_AFIADDR_bus),
	.afiba(hmc_inst_AFIBA_bus),
	.aficke(hmc_inst_AFICKE_bus),
	.aficsn(hmc_inst_AFICSN_bus),
	.afictllongidle(),
	.afictlrefreshdone(),
	.afidm(hmc_inst_AFIDM_bus),
	.afidqsburst(hmc_inst_AFIDQSBURST_bus),
	.afiodt(hmc_inst_AFIODT_bus),
	.afirdataen(hmc_inst_AFIRDATAEN_bus),
	.afirdataenfull(hmc_inst_AFIRDATAENFULL_bus),
	.afiwdata(hmc_inst_AFIWDATA_bus),
	.afiwdatavalid(hmc_inst_AFIWDATAVALID_bus),
	.bondingout1(),
	.bondingout2(),
	.bondingout3(),
	.cfgaddlat(hmc_inst_CFGADDLAT_bus),
	.cfgbankaddrwidth(hmc_inst_CFGBANKADDRWIDTH_bus),
	.cfgcaswrlat(hmc_inst_CFGCASWRLAT_bus),
	.cfgcoladdrwidth(hmc_inst_CFGCOLADDRWIDTH_bus),
	.cfgcsaddrwidth(hmc_inst_CFGCSADDRWIDTH_bus),
	.cfgdevicewidth(hmc_inst_CFGDEVICEWIDTH_bus),
	.cfginterfacewidth(hmc_inst_CFGINTERFACEWIDTH_bus),
	.cfgrowaddrwidth(hmc_inst_CFGROWADDRWIDTH_bus),
	.cfgtcl(hmc_inst_CFGTCL_bus),
	.cfgtmrd(hmc_inst_CFGTMRD_bus),
	.cfgtrefi(hmc_inst_CFGTREFI_bus),
	.cfgtrfc(hmc_inst_CFGTRFC_bus),
	.cfgtwr(hmc_inst_CFGTWR_bus),
	.ctlcalbytelaneseln(),
	.ctlmemclkdisable(hmc_inst_CTLMEMCLKDISABLE_bus),
	.dramconfig(hmc_inst_DRAMCONFIG_bus),
	.mmrrdata(),
	.ordavstdata0(),
	.ordavstdata1(),
	.ordavstdata2(),
	.ordavstdata3(),
	.scrdata());
defparam hmc_inst.attr_counter_one_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_reset = "disabled";
defparam hmc_inst.attr_counter_zero_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_reset = "disabled";
defparam hmc_inst.attr_debug_select_byte = 32'b00000000000000000000000000000000;
defparam hmc_inst.attr_static_config_valid = "disabled";
defparam hmc_inst.auto_pch_enable_0 = "disabled";
defparam hmc_inst.auto_pch_enable_1 = "disabled";
defparam hmc_inst.auto_pch_enable_2 = "disabled";
defparam hmc_inst.auto_pch_enable_3 = "disabled";
defparam hmc_inst.auto_pch_enable_4 = "disabled";
defparam hmc_inst.auto_pch_enable_5 = "disabled";
defparam hmc_inst.cal_req = "disabled";
defparam hmc_inst.cfg_burst_length = "bl_8";
defparam hmc_inst.cfg_interface_width = "dwidth_32";
defparam hmc_inst.cfg_self_rfsh_exit_cycles = "self_rfsh_exit_cycles_512";
defparam hmc_inst.cfg_starve_limit = "starve_limit_10";
defparam hmc_inst.cfg_type = "ddr3";
defparam hmc_inst.clr_intr = "no_clr_intr";
defparam hmc_inst.cmd_port_in_use_0 = "false";
defparam hmc_inst.cmd_port_in_use_1 = "false";
defparam hmc_inst.cmd_port_in_use_2 = "false";
defparam hmc_inst.cmd_port_in_use_3 = "false";
defparam hmc_inst.cmd_port_in_use_4 = "false";
defparam hmc_inst.cmd_port_in_use_5 = "false";
defparam hmc_inst.cport0_rdy_almost_full = "not_full";
defparam hmc_inst.cport0_rfifo_map = "fifo_0";
defparam hmc_inst.cport0_type = "disable";
defparam hmc_inst.cport0_wfifo_map = "fifo_0";
defparam hmc_inst.cport1_rdy_almost_full = "not_full";
defparam hmc_inst.cport1_rfifo_map = "fifo_0";
defparam hmc_inst.cport1_type = "disable";
defparam hmc_inst.cport1_wfifo_map = "fifo_0";
defparam hmc_inst.cport2_rdy_almost_full = "not_full";
defparam hmc_inst.cport2_rfifo_map = "fifo_0";
defparam hmc_inst.cport2_type = "disable";
defparam hmc_inst.cport2_wfifo_map = "fifo_0";
defparam hmc_inst.cport3_rdy_almost_full = "not_full";
defparam hmc_inst.cport3_rfifo_map = "fifo_0";
defparam hmc_inst.cport3_type = "disable";
defparam hmc_inst.cport3_wfifo_map = "fifo_0";
defparam hmc_inst.cport4_rdy_almost_full = "not_full";
defparam hmc_inst.cport4_rfifo_map = "fifo_0";
defparam hmc_inst.cport4_type = "disable";
defparam hmc_inst.cport4_wfifo_map = "fifo_0";
defparam hmc_inst.cport5_rdy_almost_full = "not_full";
defparam hmc_inst.cport5_rfifo_map = "fifo_0";
defparam hmc_inst.cport5_type = "disable";
defparam hmc_inst.cport5_wfifo_map = "fifo_0";
defparam hmc_inst.ctl_addr_order = "chip_row_bank_col";
defparam hmc_inst.ctl_ecc_enabled = "ctl_ecc_disabled";
defparam hmc_inst.ctl_ecc_rmw_enabled = "ctl_ecc_rmw_disabled";
defparam hmc_inst.ctl_regdimm_enabled = "regdimm_disabled";
defparam hmc_inst.ctl_usr_refresh = "ctl_usr_refresh_disabled";
defparam hmc_inst.ctrl_width = "data_width_64_bit";
defparam hmc_inst.cyc_to_rld_jars_0 = 1;
defparam hmc_inst.cyc_to_rld_jars_1 = 1;
defparam hmc_inst.cyc_to_rld_jars_2 = 1;
defparam hmc_inst.cyc_to_rld_jars_3 = 1;
defparam hmc_inst.cyc_to_rld_jars_4 = 1;
defparam hmc_inst.cyc_to_rld_jars_5 = 1;
defparam hmc_inst.delay_bonding = "bonding_latency_0";
defparam hmc_inst.dfx_bypass_enable = "dfx_bypass_disabled";
defparam hmc_inst.disable_merging = "merging_enabled";
defparam hmc_inst.ecc_dq_width = "ecc_dq_width_0";
defparam hmc_inst.enable_atpg = "disabled";
defparam hmc_inst.enable_bonding_0 = "disabled";
defparam hmc_inst.enable_bonding_1 = "disabled";
defparam hmc_inst.enable_bonding_2 = "disabled";
defparam hmc_inst.enable_bonding_3 = "disabled";
defparam hmc_inst.enable_bonding_4 = "disabled";
defparam hmc_inst.enable_bonding_5 = "disabled";
defparam hmc_inst.enable_bonding_wrapback = "disabled";
defparam hmc_inst.enable_burst_interrupt = "disabled";
defparam hmc_inst.enable_burst_terminate = "disabled";
defparam hmc_inst.enable_dqs_tracking = "enabled";
defparam hmc_inst.enable_ecc_code_overwrites = "disabled";
defparam hmc_inst.enable_fast_exit_ppd = "disabled";
defparam hmc_inst.enable_intr = "disabled";
defparam hmc_inst.enable_no_dm = "disabled";
defparam hmc_inst.enable_pipelineglobal = "disabled";
defparam hmc_inst.extra_ctl_clk_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_act_to_act_diff_bank = 0;
defparam hmc_inst.extra_ctl_clk_act_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_act_to_rdwr = 0;
defparam hmc_inst.extra_ctl_clk_arf_period = 0;
defparam hmc_inst.extra_ctl_clk_arf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_four_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_pch_all_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pch_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pdn_period = 0;
defparam hmc_inst.extra_ctl_clk_pdn_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd_diff_chip = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_wr = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_bc = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_diff_chip = 2;
defparam hmc_inst.extra_ctl_clk_srf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_srf_to_zq_cal = 0;
defparam hmc_inst.extra_ctl_clk_wr_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_rd = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_bc = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_diff_chip = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_wr = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_wr_diff_chip = 0;
defparam hmc_inst.gen_dbe = "gen_dbe_disabled";
defparam hmc_inst.gen_sbe = "gen_sbe_disabled";
defparam hmc_inst.inc_sync = "fifo_set_2";
defparam hmc_inst.local_if_cs_width = "addr_width_0";
defparam hmc_inst.mask_corr_dropped_intr = "disabled";
defparam hmc_inst.mask_dbe_intr = "disabled";
defparam hmc_inst.mask_sbe_intr = "disabled";
defparam hmc_inst.mem_auto_pd_cycles = 0;
defparam hmc_inst.mem_clk_entry_cycles = 10;
defparam hmc_inst.mem_if_al = "al_0";
defparam hmc_inst.mem_if_bankaddr_width = "addr_width_3";
defparam hmc_inst.mem_if_burstlength = "mem_if_burstlength_8";
defparam hmc_inst.mem_if_coladdr_width = "addr_width_10";
defparam hmc_inst.mem_if_cs_per_rank = "mem_if_cs_per_rank_1";
defparam hmc_inst.mem_if_cs_width = "mem_if_cs_width_1";
defparam hmc_inst.mem_if_dq_per_chip = "mem_if_dq_per_chip_8";
defparam hmc_inst.mem_if_dqs_width = "dqs_width_4";
defparam hmc_inst.mem_if_dwidth = "mem_if_dwidth_32";
defparam hmc_inst.mem_if_memtype = "ddr3_sdram";
defparam hmc_inst.mem_if_rowaddr_width = "addr_width_15";
defparam hmc_inst.mem_if_speedbin = "ddr3_1600_8_8_8";
defparam hmc_inst.mem_if_tccd = "tccd_4";
defparam hmc_inst.mem_if_tcl = "tcl_11";
defparam hmc_inst.mem_if_tcwl = "tcwl_8";
defparam hmc_inst.mem_if_tfaw = "tfaw_12";
defparam hmc_inst.mem_if_tmrd = "tmrd_4";
defparam hmc_inst.mem_if_tras = "tras_14";
defparam hmc_inst.mem_if_trc = "trc_20";
defparam hmc_inst.mem_if_trcd = "trcd_6";
defparam hmc_inst.mem_if_trefi = 3120;
defparam hmc_inst.mem_if_trfc = 104;
defparam hmc_inst.mem_if_trp = "trp_6";
defparam hmc_inst.mem_if_trrd = "trrd_3";
defparam hmc_inst.mem_if_trtp = "trtp_3";
defparam hmc_inst.mem_if_twr = "twr_6";
defparam hmc_inst.mem_if_twtr = "twtr_4";
defparam hmc_inst.mmr_cfg_mem_bl = "mp_bl_8";
defparam hmc_inst.output_regd = "disabled";
defparam hmc_inst.pdn_exit_cycles = "slow_exit";
defparam hmc_inst.port0_width = "port_32_bit";
defparam hmc_inst.port1_width = "port_32_bit";
defparam hmc_inst.port2_width = "port_32_bit";
defparam hmc_inst.port3_width = "port_32_bit";
defparam hmc_inst.port4_width = "port_32_bit";
defparam hmc_inst.port5_width = "port_32_bit";
defparam hmc_inst.power_saving_exit_cycles = 5;
defparam hmc_inst.priority_0_0 = "weight_0";
defparam hmc_inst.priority_0_1 = "weight_0";
defparam hmc_inst.priority_0_2 = "weight_0";
defparam hmc_inst.priority_0_3 = "weight_0";
defparam hmc_inst.priority_0_4 = "weight_0";
defparam hmc_inst.priority_0_5 = "weight_0";
defparam hmc_inst.priority_1_0 = "weight_0";
defparam hmc_inst.priority_1_1 = "weight_0";
defparam hmc_inst.priority_1_2 = "weight_0";
defparam hmc_inst.priority_1_3 = "weight_0";
defparam hmc_inst.priority_1_4 = "weight_0";
defparam hmc_inst.priority_1_5 = "weight_0";
defparam hmc_inst.priority_2_0 = "weight_0";
defparam hmc_inst.priority_2_1 = "weight_0";
defparam hmc_inst.priority_2_2 = "weight_0";
defparam hmc_inst.priority_2_3 = "weight_0";
defparam hmc_inst.priority_2_4 = "weight_0";
defparam hmc_inst.priority_2_5 = "weight_0";
defparam hmc_inst.priority_3_0 = "weight_0";
defparam hmc_inst.priority_3_1 = "weight_0";
defparam hmc_inst.priority_3_2 = "weight_0";
defparam hmc_inst.priority_3_3 = "weight_0";
defparam hmc_inst.priority_3_4 = "weight_0";
defparam hmc_inst.priority_3_5 = "weight_0";
defparam hmc_inst.priority_4_0 = "weight_0";
defparam hmc_inst.priority_4_1 = "weight_0";
defparam hmc_inst.priority_4_2 = "weight_0";
defparam hmc_inst.priority_4_3 = "weight_0";
defparam hmc_inst.priority_4_4 = "weight_0";
defparam hmc_inst.priority_4_5 = "weight_0";
defparam hmc_inst.priority_5_0 = "weight_0";
defparam hmc_inst.priority_5_1 = "weight_0";
defparam hmc_inst.priority_5_2 = "weight_0";
defparam hmc_inst.priority_5_3 = "weight_0";
defparam hmc_inst.priority_5_4 = "weight_0";
defparam hmc_inst.priority_5_5 = "weight_0";
defparam hmc_inst.priority_6_0 = "weight_0";
defparam hmc_inst.priority_6_1 = "weight_0";
defparam hmc_inst.priority_6_2 = "weight_0";
defparam hmc_inst.priority_6_3 = "weight_0";
defparam hmc_inst.priority_6_4 = "weight_0";
defparam hmc_inst.priority_6_5 = "weight_0";
defparam hmc_inst.priority_7_0 = "weight_0";
defparam hmc_inst.priority_7_1 = "weight_0";
defparam hmc_inst.priority_7_2 = "weight_0";
defparam hmc_inst.priority_7_3 = "weight_0";
defparam hmc_inst.priority_7_4 = "weight_0";
defparam hmc_inst.priority_7_5 = "weight_0";
defparam hmc_inst.priority_remap = 0;
defparam hmc_inst.rcfg_static_weight_0 = "weight_0";
defparam hmc_inst.rcfg_static_weight_1 = "weight_0";
defparam hmc_inst.rcfg_static_weight_2 = "weight_0";
defparam hmc_inst.rcfg_static_weight_3 = "weight_0";
defparam hmc_inst.rcfg_static_weight_4 = "weight_0";
defparam hmc_inst.rcfg_static_weight_5 = "weight_0";
defparam hmc_inst.rcfg_sum_wt_priority_0 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_1 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_2 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_3 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_4 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_5 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_6 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_7 = 0;
defparam hmc_inst.rcfg_user_priority_0 = "priority_1";
defparam hmc_inst.rcfg_user_priority_1 = "priority_1";
defparam hmc_inst.rcfg_user_priority_2 = "priority_1";
defparam hmc_inst.rcfg_user_priority_3 = "priority_1";
defparam hmc_inst.rcfg_user_priority_4 = "priority_1";
defparam hmc_inst.rcfg_user_priority_5 = "priority_1";
defparam hmc_inst.rd_dwidth_0 = "dwidth_0";
defparam hmc_inst.rd_dwidth_1 = "dwidth_0";
defparam hmc_inst.rd_dwidth_2 = "dwidth_0";
defparam hmc_inst.rd_dwidth_3 = "dwidth_0";
defparam hmc_inst.rd_dwidth_4 = "dwidth_0";
defparam hmc_inst.rd_dwidth_5 = "dwidth_0";
defparam hmc_inst.rd_fifo_in_use_0 = "false";
defparam hmc_inst.rd_fifo_in_use_1 = "false";
defparam hmc_inst.rd_fifo_in_use_2 = "false";
defparam hmc_inst.rd_fifo_in_use_3 = "false";
defparam hmc_inst.rd_port_info_0 = "use_no";
defparam hmc_inst.rd_port_info_1 = "use_no";
defparam hmc_inst.rd_port_info_2 = "use_no";
defparam hmc_inst.rd_port_info_3 = "use_no";
defparam hmc_inst.rd_port_info_4 = "use_no";
defparam hmc_inst.rd_port_info_5 = "use_no";
defparam hmc_inst.read_odt_chip = "odt_disabled";
defparam hmc_inst.reorder_data = "data_reordering";
defparam hmc_inst.rfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.single_ready_0 = "concatenate_rdy";
defparam hmc_inst.single_ready_1 = "concatenate_rdy";
defparam hmc_inst.single_ready_2 = "concatenate_rdy";
defparam hmc_inst.single_ready_3 = "concatenate_rdy";
defparam hmc_inst.static_weight_0 = "weight_0";
defparam hmc_inst.static_weight_1 = "weight_0";
defparam hmc_inst.static_weight_2 = "weight_0";
defparam hmc_inst.static_weight_3 = "weight_0";
defparam hmc_inst.static_weight_4 = "weight_0";
defparam hmc_inst.static_weight_5 = "weight_0";
defparam hmc_inst.sum_wt_priority_0 = 0;
defparam hmc_inst.sum_wt_priority_1 = 0;
defparam hmc_inst.sum_wt_priority_2 = 0;
defparam hmc_inst.sum_wt_priority_3 = 0;
defparam hmc_inst.sum_wt_priority_4 = 0;
defparam hmc_inst.sum_wt_priority_5 = 0;
defparam hmc_inst.sum_wt_priority_6 = 0;
defparam hmc_inst.sum_wt_priority_7 = 0;
defparam hmc_inst.sync_mode_0 = "asynchronous";
defparam hmc_inst.sync_mode_1 = "asynchronous";
defparam hmc_inst.sync_mode_2 = "asynchronous";
defparam hmc_inst.sync_mode_3 = "asynchronous";
defparam hmc_inst.sync_mode_4 = "asynchronous";
defparam hmc_inst.sync_mode_5 = "asynchronous";
defparam hmc_inst.test_mode = "normal_mode";
defparam hmc_inst.thld_jar1_0 = "threshold_32";
defparam hmc_inst.thld_jar1_1 = "threshold_32";
defparam hmc_inst.thld_jar1_2 = "threshold_32";
defparam hmc_inst.thld_jar1_3 = "threshold_32";
defparam hmc_inst.thld_jar1_4 = "threshold_32";
defparam hmc_inst.thld_jar1_5 = "threshold_32";
defparam hmc_inst.thld_jar2_0 = "threshold_16";
defparam hmc_inst.thld_jar2_1 = "threshold_16";
defparam hmc_inst.thld_jar2_2 = "threshold_16";
defparam hmc_inst.thld_jar2_3 = "threshold_16";
defparam hmc_inst.thld_jar2_4 = "threshold_16";
defparam hmc_inst.thld_jar2_5 = "threshold_16";
defparam hmc_inst.use_almost_empty_0 = "empty";
defparam hmc_inst.use_almost_empty_1 = "empty";
defparam hmc_inst.use_almost_empty_2 = "empty";
defparam hmc_inst.use_almost_empty_3 = "empty";
defparam hmc_inst.user_ecc_en = "disable";
defparam hmc_inst.user_priority_0 = "priority_1";
defparam hmc_inst.user_priority_1 = "priority_1";
defparam hmc_inst.user_priority_2 = "priority_1";
defparam hmc_inst.user_priority_3 = "priority_1";
defparam hmc_inst.user_priority_4 = "priority_1";
defparam hmc_inst.user_priority_5 = "priority_1";
defparam hmc_inst.wfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo0_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo1_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo2_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo3_rdy_almost_full = "not_full";
defparam hmc_inst.wr_dwidth_0 = "dwidth_0";
defparam hmc_inst.wr_dwidth_1 = "dwidth_0";
defparam hmc_inst.wr_dwidth_2 = "dwidth_0";
defparam hmc_inst.wr_dwidth_3 = "dwidth_0";
defparam hmc_inst.wr_dwidth_4 = "dwidth_0";
defparam hmc_inst.wr_dwidth_5 = "dwidth_0";
defparam hmc_inst.wr_fifo_in_use_0 = "false";
defparam hmc_inst.wr_fifo_in_use_1 = "false";
defparam hmc_inst.wr_fifo_in_use_2 = "false";
defparam hmc_inst.wr_fifo_in_use_3 = "false";
defparam hmc_inst.wr_port_info_0 = "use_no";
defparam hmc_inst.wr_port_info_1 = "use_no";
defparam hmc_inst.wr_port_info_2 = "use_no";
defparam hmc_inst.wr_port_info_3 = "use_no";
defparam hmc_inst.wr_port_info_4 = "use_no";
defparam hmc_inst.wr_port_info_5 = "use_no";
defparam hmc_inst.write_odt_chip = "write_chip0_odt0_chip1";

endmodule

module Computer_System_altera_mem_if_oct_cyclonev (
	parallelterminationcontrol,
	seriesterminationcontrol,
	oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[15:0] parallelterminationcontrol;
output 	[15:0] seriesterminationcontrol;
input 	oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sd1a_0~O_CLKUSRDFTOUT ;
wire \wire_sd1a_serdataout[0] ;

wire [15:0] sd2a_0_PARALLELTERMINATIONCONTROL_bus;
wire [15:0] sd2a_0_SERIESTERMINATIONCONTROL_bus;

assign parallelterminationcontrol[0] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[0];
assign parallelterminationcontrol[1] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[1];
assign parallelterminationcontrol[2] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[2];
assign parallelterminationcontrol[3] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[3];
assign parallelterminationcontrol[4] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[4];
assign parallelterminationcontrol[5] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[5];
assign parallelterminationcontrol[6] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[6];
assign parallelterminationcontrol[7] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[7];
assign parallelterminationcontrol[8] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[8];
assign parallelterminationcontrol[9] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[9];
assign parallelterminationcontrol[10] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[10];
assign parallelterminationcontrol[11] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[11];
assign parallelterminationcontrol[12] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[12];
assign parallelterminationcontrol[13] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[13];
assign parallelterminationcontrol[14] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[14];
assign parallelterminationcontrol[15] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[15];

assign seriesterminationcontrol[0] = sd2a_0_SERIESTERMINATIONCONTROL_bus[0];
assign seriesterminationcontrol[1] = sd2a_0_SERIESTERMINATIONCONTROL_bus[1];
assign seriesterminationcontrol[2] = sd2a_0_SERIESTERMINATIONCONTROL_bus[2];
assign seriesterminationcontrol[3] = sd2a_0_SERIESTERMINATIONCONTROL_bus[3];
assign seriesterminationcontrol[4] = sd2a_0_SERIESTERMINATIONCONTROL_bus[4];
assign seriesterminationcontrol[5] = sd2a_0_SERIESTERMINATIONCONTROL_bus[5];
assign seriesterminationcontrol[6] = sd2a_0_SERIESTERMINATIONCONTROL_bus[6];
assign seriesterminationcontrol[7] = sd2a_0_SERIESTERMINATIONCONTROL_bus[7];
assign seriesterminationcontrol[8] = sd2a_0_SERIESTERMINATIONCONTROL_bus[8];
assign seriesterminationcontrol[9] = sd2a_0_SERIESTERMINATIONCONTROL_bus[9];
assign seriesterminationcontrol[10] = sd2a_0_SERIESTERMINATIONCONTROL_bus[10];
assign seriesterminationcontrol[11] = sd2a_0_SERIESTERMINATIONCONTROL_bus[11];
assign seriesterminationcontrol[12] = sd2a_0_SERIESTERMINATIONCONTROL_bus[12];
assign seriesterminationcontrol[13] = sd2a_0_SERIESTERMINATIONCONTROL_bus[13];
assign seriesterminationcontrol[14] = sd2a_0_SERIESTERMINATIONCONTROL_bus[14];
assign seriesterminationcontrol[15] = sd2a_0_SERIESTERMINATIONCONTROL_bus[15];

cyclonev_termination_logic sd2a_0(
	.s2pload(gnd),
	.scanclk(gnd),
	.scanenable(gnd),
	.serdata(\wire_sd1a_serdataout[0] ),
	.enser(4'b0000),
	.parallelterminationcontrol(sd2a_0_PARALLELTERMINATIONCONTROL_bus),
	.seriesterminationcontrol(sd2a_0_SERIESTERMINATIONCONTROL_bus));

cyclonev_termination sd1a_0(
	.clkenusr(gnd),
	.clkusr(gnd),
	.enserusr(gnd),
	.nclrusr(gnd),
	.rzqin(oct_rzqin),
	.scanclk(gnd),
	.scanen(gnd),
	.scanin(gnd),
	.serdatafromcore(gnd),
	.serdatain(gnd),
	.otherenser(10'b0000000000),
	.clkusrdftout(\sd1a_0~O_CLKUSRDFTOUT ),
	.compoutrdn(),
	.compoutrup(),
	.enserout(),
	.scanout(),
	.serdataout(\wire_sd1a_serdataout[0] ),
	.serdatatocore());

endmodule

module Computer_System_hps_sdram_p0 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid_0,
	ctl_reset_n,
	afi_rdata_0,
	afi_rdata_1,
	afi_rdata_2,
	afi_rdata_3,
	afi_rdata_4,
	afi_rdata_5,
	afi_rdata_6,
	afi_rdata_7,
	afi_rdata_8,
	afi_rdata_9,
	afi_rdata_10,
	afi_rdata_11,
	afi_rdata_12,
	afi_rdata_13,
	afi_rdata_14,
	afi_rdata_15,
	afi_rdata_16,
	afi_rdata_17,
	afi_rdata_18,
	afi_rdata_19,
	afi_rdata_20,
	afi_rdata_21,
	afi_rdata_22,
	afi_rdata_23,
	afi_rdata_24,
	afi_rdata_25,
	afi_rdata_26,
	afi_rdata_27,
	afi_rdata_28,
	afi_rdata_29,
	afi_rdata_30,
	afi_rdata_31,
	afi_rdata_32,
	afi_rdata_33,
	afi_rdata_34,
	afi_rdata_35,
	afi_rdata_36,
	afi_rdata_37,
	afi_rdata_38,
	afi_rdata_39,
	afi_rdata_40,
	afi_rdata_41,
	afi_rdata_42,
	afi_rdata_43,
	afi_rdata_44,
	afi_rdata_45,
	afi_rdata_46,
	afi_rdata_47,
	afi_rdata_48,
	afi_rdata_49,
	afi_rdata_50,
	afi_rdata_51,
	afi_rdata_52,
	afi_rdata_53,
	afi_rdata_54,
	afi_rdata_55,
	afi_rdata_56,
	afi_rdata_57,
	afi_rdata_58,
	afi_rdata_59,
	afi_rdata_60,
	afi_rdata_61,
	afi_rdata_62,
	afi_rdata_63,
	afi_rdata_64,
	afi_rdata_65,
	afi_rdata_66,
	afi_rdata_67,
	afi_rdata_68,
	afi_rdata_69,
	afi_rdata_70,
	afi_rdata_71,
	afi_rdata_72,
	afi_rdata_73,
	afi_rdata_74,
	afi_rdata_75,
	afi_rdata_76,
	afi_rdata_77,
	afi_rdata_78,
	afi_rdata_79,
	afi_wlat_0,
	afi_wlat_1,
	afi_wlat_2,
	afi_wlat_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n_0,
	afi_ras_n_0,
	afi_rst_n_0,
	afi_we_n_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_addr_14,
	afi_addr_15,
	afi_addr_16,
	afi_addr_17,
	afi_addr_18,
	afi_addr_19,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_cke_0,
	afi_cke_1,
	afi_cs_n_0,
	afi_cs_n_1,
	afi_dm_int_0,
	afi_dm_int_1,
	afi_dm_int_2,
	afi_dm_int_3,
	afi_dm_int_4,
	afi_dm_int_5,
	afi_dm_int_6,
	afi_dm_int_7,
	afi_dm_int_8,
	afi_dm_int_9,
	afi_dqs_burst_0,
	afi_dqs_burst_1,
	afi_dqs_burst_2,
	afi_dqs_burst_3,
	afi_dqs_burst_4,
	afi_odt_0,
	afi_odt_1,
	afi_rdata_en_0,
	afi_rdata_en_1,
	afi_rdata_en_2,
	afi_rdata_en_3,
	afi_rdata_en_4,
	afi_rdata_en_full_0,
	afi_rdata_en_full_1,
	afi_rdata_en_full_2,
	afi_rdata_en_full_3,
	afi_rdata_en_full_4,
	afi_wdata_int_0,
	afi_wdata_int_1,
	afi_wdata_int_2,
	afi_wdata_int_3,
	afi_wdata_int_4,
	afi_wdata_int_5,
	afi_wdata_int_6,
	afi_wdata_int_7,
	afi_wdata_int_8,
	afi_wdata_int_9,
	afi_wdata_int_10,
	afi_wdata_int_11,
	afi_wdata_int_12,
	afi_wdata_int_13,
	afi_wdata_int_14,
	afi_wdata_int_15,
	afi_wdata_int_16,
	afi_wdata_int_17,
	afi_wdata_int_18,
	afi_wdata_int_19,
	afi_wdata_int_20,
	afi_wdata_int_21,
	afi_wdata_int_22,
	afi_wdata_int_23,
	afi_wdata_int_24,
	afi_wdata_int_25,
	afi_wdata_int_26,
	afi_wdata_int_27,
	afi_wdata_int_28,
	afi_wdata_int_29,
	afi_wdata_int_30,
	afi_wdata_int_31,
	afi_wdata_int_32,
	afi_wdata_int_33,
	afi_wdata_int_34,
	afi_wdata_int_35,
	afi_wdata_int_36,
	afi_wdata_int_37,
	afi_wdata_int_38,
	afi_wdata_int_39,
	afi_wdata_int_40,
	afi_wdata_int_41,
	afi_wdata_int_42,
	afi_wdata_int_43,
	afi_wdata_int_44,
	afi_wdata_int_45,
	afi_wdata_int_46,
	afi_wdata_int_47,
	afi_wdata_int_48,
	afi_wdata_int_49,
	afi_wdata_int_50,
	afi_wdata_int_51,
	afi_wdata_int_52,
	afi_wdata_int_53,
	afi_wdata_int_54,
	afi_wdata_int_55,
	afi_wdata_int_56,
	afi_wdata_int_57,
	afi_wdata_int_58,
	afi_wdata_int_59,
	afi_wdata_int_60,
	afi_wdata_int_61,
	afi_wdata_int_62,
	afi_wdata_int_63,
	afi_wdata_int_64,
	afi_wdata_int_65,
	afi_wdata_int_66,
	afi_wdata_int_67,
	afi_wdata_int_68,
	afi_wdata_int_69,
	afi_wdata_int_70,
	afi_wdata_int_71,
	afi_wdata_int_72,
	afi_wdata_int_73,
	afi_wdata_int_74,
	afi_wdata_int_75,
	afi_wdata_int_76,
	afi_wdata_int_77,
	afi_wdata_int_78,
	afi_wdata_int_79,
	afi_wdata_valid_0,
	afi_wdata_valid_1,
	afi_wdata_valid_2,
	afi_wdata_valid_3,
	afi_wdata_valid_4,
	cfg_addlat_wire_0,
	cfg_addlat_wire_1,
	cfg_addlat_wire_2,
	cfg_addlat_wire_3,
	cfg_addlat_wire_4,
	cfg_bankaddrwidth_wire_0,
	cfg_bankaddrwidth_wire_1,
	cfg_bankaddrwidth_wire_2,
	cfg_caswrlat_wire_0,
	cfg_caswrlat_wire_1,
	cfg_caswrlat_wire_2,
	cfg_caswrlat_wire_3,
	cfg_coladdrwidth_wire_0,
	cfg_coladdrwidth_wire_1,
	cfg_coladdrwidth_wire_2,
	cfg_coladdrwidth_wire_3,
	cfg_coladdrwidth_wire_4,
	cfg_csaddrwidth_wire_0,
	cfg_csaddrwidth_wire_1,
	cfg_csaddrwidth_wire_2,
	cfg_devicewidth_wire_0,
	cfg_devicewidth_wire_1,
	cfg_devicewidth_wire_2,
	cfg_devicewidth_wire_3,
	cfg_interfacewidth_wire_0,
	cfg_interfacewidth_wire_1,
	cfg_interfacewidth_wire_2,
	cfg_interfacewidth_wire_3,
	cfg_interfacewidth_wire_4,
	cfg_interfacewidth_wire_5,
	cfg_interfacewidth_wire_6,
	cfg_interfacewidth_wire_7,
	cfg_rowaddrwidth_wire_0,
	cfg_rowaddrwidth_wire_1,
	cfg_rowaddrwidth_wire_2,
	cfg_rowaddrwidth_wire_3,
	cfg_rowaddrwidth_wire_4,
	cfg_tcl_wire_0,
	cfg_tcl_wire_1,
	cfg_tcl_wire_2,
	cfg_tcl_wire_3,
	cfg_tcl_wire_4,
	cfg_tmrd_wire_0,
	cfg_tmrd_wire_1,
	cfg_tmrd_wire_2,
	cfg_tmrd_wire_3,
	cfg_trefi_wire_0,
	cfg_trefi_wire_1,
	cfg_trefi_wire_2,
	cfg_trefi_wire_3,
	cfg_trefi_wire_4,
	cfg_trefi_wire_5,
	cfg_trefi_wire_6,
	cfg_trefi_wire_7,
	cfg_trefi_wire_8,
	cfg_trefi_wire_9,
	cfg_trefi_wire_10,
	cfg_trefi_wire_11,
	cfg_trefi_wire_12,
	cfg_trfc_wire_0,
	cfg_trfc_wire_1,
	cfg_trfc_wire_2,
	cfg_trfc_wire_3,
	cfg_trfc_wire_4,
	cfg_trfc_wire_5,
	cfg_trfc_wire_6,
	cfg_trfc_wire_7,
	cfg_twr_wire_0,
	cfg_twr_wire_1,
	cfg_twr_wire_2,
	cfg_twr_wire_3,
	afi_mem_clk_disable_0,
	cfg_dramconfig_wire_0,
	cfg_dramconfig_wire_1,
	cfg_dramconfig_wire_2,
	cfg_dramconfig_wire_3,
	cfg_dramconfig_wire_4,
	cfg_dramconfig_wire_5,
	cfg_dramconfig_wire_6,
	cfg_dramconfig_wire_7,
	cfg_dramconfig_wire_8,
	cfg_dramconfig_wire_9,
	cfg_dramconfig_wire_10,
	cfg_dramconfig_wire_11,
	cfg_dramconfig_wire_12,
	cfg_dramconfig_wire_13,
	cfg_dramconfig_wire_14,
	cfg_dramconfig_wire_15,
	cfg_dramconfig_wire_16,
	cfg_dramconfig_wire_17,
	cfg_dramconfig_wire_18,
	cfg_dramconfig_wire_19,
	cfg_dramconfig_wire_20,
	ctl_clk,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	afi_rdata_valid_0;
output 	ctl_reset_n;
output 	afi_rdata_0;
output 	afi_rdata_1;
output 	afi_rdata_2;
output 	afi_rdata_3;
output 	afi_rdata_4;
output 	afi_rdata_5;
output 	afi_rdata_6;
output 	afi_rdata_7;
output 	afi_rdata_8;
output 	afi_rdata_9;
output 	afi_rdata_10;
output 	afi_rdata_11;
output 	afi_rdata_12;
output 	afi_rdata_13;
output 	afi_rdata_14;
output 	afi_rdata_15;
output 	afi_rdata_16;
output 	afi_rdata_17;
output 	afi_rdata_18;
output 	afi_rdata_19;
output 	afi_rdata_20;
output 	afi_rdata_21;
output 	afi_rdata_22;
output 	afi_rdata_23;
output 	afi_rdata_24;
output 	afi_rdata_25;
output 	afi_rdata_26;
output 	afi_rdata_27;
output 	afi_rdata_28;
output 	afi_rdata_29;
output 	afi_rdata_30;
output 	afi_rdata_31;
output 	afi_rdata_32;
output 	afi_rdata_33;
output 	afi_rdata_34;
output 	afi_rdata_35;
output 	afi_rdata_36;
output 	afi_rdata_37;
output 	afi_rdata_38;
output 	afi_rdata_39;
output 	afi_rdata_40;
output 	afi_rdata_41;
output 	afi_rdata_42;
output 	afi_rdata_43;
output 	afi_rdata_44;
output 	afi_rdata_45;
output 	afi_rdata_46;
output 	afi_rdata_47;
output 	afi_rdata_48;
output 	afi_rdata_49;
output 	afi_rdata_50;
output 	afi_rdata_51;
output 	afi_rdata_52;
output 	afi_rdata_53;
output 	afi_rdata_54;
output 	afi_rdata_55;
output 	afi_rdata_56;
output 	afi_rdata_57;
output 	afi_rdata_58;
output 	afi_rdata_59;
output 	afi_rdata_60;
output 	afi_rdata_61;
output 	afi_rdata_62;
output 	afi_rdata_63;
output 	afi_rdata_64;
output 	afi_rdata_65;
output 	afi_rdata_66;
output 	afi_rdata_67;
output 	afi_rdata_68;
output 	afi_rdata_69;
output 	afi_rdata_70;
output 	afi_rdata_71;
output 	afi_rdata_72;
output 	afi_rdata_73;
output 	afi_rdata_74;
output 	afi_rdata_75;
output 	afi_rdata_76;
output 	afi_rdata_77;
output 	afi_rdata_78;
output 	afi_rdata_79;
output 	afi_wlat_0;
output 	afi_wlat_1;
output 	afi_wlat_2;
output 	afi_wlat_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	afi_cas_n_0;
input 	afi_ras_n_0;
input 	afi_rst_n_0;
input 	afi_we_n_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_addr_14;
input 	afi_addr_15;
input 	afi_addr_16;
input 	afi_addr_17;
input 	afi_addr_18;
input 	afi_addr_19;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_cke_0;
input 	afi_cke_1;
input 	afi_cs_n_0;
input 	afi_cs_n_1;
input 	afi_dm_int_0;
input 	afi_dm_int_1;
input 	afi_dm_int_2;
input 	afi_dm_int_3;
input 	afi_dm_int_4;
input 	afi_dm_int_5;
input 	afi_dm_int_6;
input 	afi_dm_int_7;
input 	afi_dm_int_8;
input 	afi_dm_int_9;
input 	afi_dqs_burst_0;
input 	afi_dqs_burst_1;
input 	afi_dqs_burst_2;
input 	afi_dqs_burst_3;
input 	afi_dqs_burst_4;
input 	afi_odt_0;
input 	afi_odt_1;
input 	afi_rdata_en_0;
input 	afi_rdata_en_1;
input 	afi_rdata_en_2;
input 	afi_rdata_en_3;
input 	afi_rdata_en_4;
input 	afi_rdata_en_full_0;
input 	afi_rdata_en_full_1;
input 	afi_rdata_en_full_2;
input 	afi_rdata_en_full_3;
input 	afi_rdata_en_full_4;
input 	afi_wdata_int_0;
input 	afi_wdata_int_1;
input 	afi_wdata_int_2;
input 	afi_wdata_int_3;
input 	afi_wdata_int_4;
input 	afi_wdata_int_5;
input 	afi_wdata_int_6;
input 	afi_wdata_int_7;
input 	afi_wdata_int_8;
input 	afi_wdata_int_9;
input 	afi_wdata_int_10;
input 	afi_wdata_int_11;
input 	afi_wdata_int_12;
input 	afi_wdata_int_13;
input 	afi_wdata_int_14;
input 	afi_wdata_int_15;
input 	afi_wdata_int_16;
input 	afi_wdata_int_17;
input 	afi_wdata_int_18;
input 	afi_wdata_int_19;
input 	afi_wdata_int_20;
input 	afi_wdata_int_21;
input 	afi_wdata_int_22;
input 	afi_wdata_int_23;
input 	afi_wdata_int_24;
input 	afi_wdata_int_25;
input 	afi_wdata_int_26;
input 	afi_wdata_int_27;
input 	afi_wdata_int_28;
input 	afi_wdata_int_29;
input 	afi_wdata_int_30;
input 	afi_wdata_int_31;
input 	afi_wdata_int_32;
input 	afi_wdata_int_33;
input 	afi_wdata_int_34;
input 	afi_wdata_int_35;
input 	afi_wdata_int_36;
input 	afi_wdata_int_37;
input 	afi_wdata_int_38;
input 	afi_wdata_int_39;
input 	afi_wdata_int_40;
input 	afi_wdata_int_41;
input 	afi_wdata_int_42;
input 	afi_wdata_int_43;
input 	afi_wdata_int_44;
input 	afi_wdata_int_45;
input 	afi_wdata_int_46;
input 	afi_wdata_int_47;
input 	afi_wdata_int_48;
input 	afi_wdata_int_49;
input 	afi_wdata_int_50;
input 	afi_wdata_int_51;
input 	afi_wdata_int_52;
input 	afi_wdata_int_53;
input 	afi_wdata_int_54;
input 	afi_wdata_int_55;
input 	afi_wdata_int_56;
input 	afi_wdata_int_57;
input 	afi_wdata_int_58;
input 	afi_wdata_int_59;
input 	afi_wdata_int_60;
input 	afi_wdata_int_61;
input 	afi_wdata_int_62;
input 	afi_wdata_int_63;
input 	afi_wdata_int_64;
input 	afi_wdata_int_65;
input 	afi_wdata_int_66;
input 	afi_wdata_int_67;
input 	afi_wdata_int_68;
input 	afi_wdata_int_69;
input 	afi_wdata_int_70;
input 	afi_wdata_int_71;
input 	afi_wdata_int_72;
input 	afi_wdata_int_73;
input 	afi_wdata_int_74;
input 	afi_wdata_int_75;
input 	afi_wdata_int_76;
input 	afi_wdata_int_77;
input 	afi_wdata_int_78;
input 	afi_wdata_int_79;
input 	afi_wdata_valid_0;
input 	afi_wdata_valid_1;
input 	afi_wdata_valid_2;
input 	afi_wdata_valid_3;
input 	afi_wdata_valid_4;
input 	cfg_addlat_wire_0;
input 	cfg_addlat_wire_1;
input 	cfg_addlat_wire_2;
input 	cfg_addlat_wire_3;
input 	cfg_addlat_wire_4;
input 	cfg_bankaddrwidth_wire_0;
input 	cfg_bankaddrwidth_wire_1;
input 	cfg_bankaddrwidth_wire_2;
input 	cfg_caswrlat_wire_0;
input 	cfg_caswrlat_wire_1;
input 	cfg_caswrlat_wire_2;
input 	cfg_caswrlat_wire_3;
input 	cfg_coladdrwidth_wire_0;
input 	cfg_coladdrwidth_wire_1;
input 	cfg_coladdrwidth_wire_2;
input 	cfg_coladdrwidth_wire_3;
input 	cfg_coladdrwidth_wire_4;
input 	cfg_csaddrwidth_wire_0;
input 	cfg_csaddrwidth_wire_1;
input 	cfg_csaddrwidth_wire_2;
input 	cfg_devicewidth_wire_0;
input 	cfg_devicewidth_wire_1;
input 	cfg_devicewidth_wire_2;
input 	cfg_devicewidth_wire_3;
input 	cfg_interfacewidth_wire_0;
input 	cfg_interfacewidth_wire_1;
input 	cfg_interfacewidth_wire_2;
input 	cfg_interfacewidth_wire_3;
input 	cfg_interfacewidth_wire_4;
input 	cfg_interfacewidth_wire_5;
input 	cfg_interfacewidth_wire_6;
input 	cfg_interfacewidth_wire_7;
input 	cfg_rowaddrwidth_wire_0;
input 	cfg_rowaddrwidth_wire_1;
input 	cfg_rowaddrwidth_wire_2;
input 	cfg_rowaddrwidth_wire_3;
input 	cfg_rowaddrwidth_wire_4;
input 	cfg_tcl_wire_0;
input 	cfg_tcl_wire_1;
input 	cfg_tcl_wire_2;
input 	cfg_tcl_wire_3;
input 	cfg_tcl_wire_4;
input 	cfg_tmrd_wire_0;
input 	cfg_tmrd_wire_1;
input 	cfg_tmrd_wire_2;
input 	cfg_tmrd_wire_3;
input 	cfg_trefi_wire_0;
input 	cfg_trefi_wire_1;
input 	cfg_trefi_wire_2;
input 	cfg_trefi_wire_3;
input 	cfg_trefi_wire_4;
input 	cfg_trefi_wire_5;
input 	cfg_trefi_wire_6;
input 	cfg_trefi_wire_7;
input 	cfg_trefi_wire_8;
input 	cfg_trefi_wire_9;
input 	cfg_trefi_wire_10;
input 	cfg_trefi_wire_11;
input 	cfg_trefi_wire_12;
input 	cfg_trfc_wire_0;
input 	cfg_trfc_wire_1;
input 	cfg_trfc_wire_2;
input 	cfg_trfc_wire_3;
input 	cfg_trfc_wire_4;
input 	cfg_trfc_wire_5;
input 	cfg_trfc_wire_6;
input 	cfg_trfc_wire_7;
input 	cfg_twr_wire_0;
input 	cfg_twr_wire_1;
input 	cfg_twr_wire_2;
input 	cfg_twr_wire_3;
input 	afi_mem_clk_disable_0;
input 	cfg_dramconfig_wire_0;
input 	cfg_dramconfig_wire_1;
input 	cfg_dramconfig_wire_2;
input 	cfg_dramconfig_wire_3;
input 	cfg_dramconfig_wire_4;
input 	cfg_dramconfig_wire_5;
input 	cfg_dramconfig_wire_6;
input 	cfg_dramconfig_wire_7;
input 	cfg_dramconfig_wire_8;
input 	cfg_dramconfig_wire_9;
input 	cfg_dramconfig_wire_10;
input 	cfg_dramconfig_wire_11;
input 	cfg_dramconfig_wire_12;
input 	cfg_dramconfig_wire_13;
input 	cfg_dramconfig_wire_14;
input 	cfg_dramconfig_wire_15;
input 	cfg_dramconfig_wire_16;
input 	cfg_dramconfig_wire_17;
input 	cfg_dramconfig_wire_18;
input 	cfg_dramconfig_wire_19;
input 	cfg_dramconfig_wire_20;
output 	ctl_clk;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_hps_sdram_p0_acv_hard_memphy umemphy(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(afi_cal_fail),
	.afi_cal_success(afi_cal_success),
	.afi_rdata_valid({afi_rdata_valid_0}),
	.ctl_reset_n(ctl_reset_n),
	.afi_rdata({afi_rdata_79,afi_rdata_78,afi_rdata_77,afi_rdata_76,afi_rdata_75,afi_rdata_74,afi_rdata_73,afi_rdata_72,afi_rdata_71,afi_rdata_70,afi_rdata_69,afi_rdata_68,afi_rdata_67,afi_rdata_66,afi_rdata_65,afi_rdata_64,afi_rdata_63,afi_rdata_62,afi_rdata_61,afi_rdata_60,afi_rdata_59,
afi_rdata_58,afi_rdata_57,afi_rdata_56,afi_rdata_55,afi_rdata_54,afi_rdata_53,afi_rdata_52,afi_rdata_51,afi_rdata_50,afi_rdata_49,afi_rdata_48,afi_rdata_47,afi_rdata_46,afi_rdata_45,afi_rdata_44,afi_rdata_43,afi_rdata_42,afi_rdata_41,afi_rdata_40,afi_rdata_39,afi_rdata_38,
afi_rdata_37,afi_rdata_36,afi_rdata_35,afi_rdata_34,afi_rdata_33,afi_rdata_32,afi_rdata_31,afi_rdata_30,afi_rdata_29,afi_rdata_28,afi_rdata_27,afi_rdata_26,afi_rdata_25,afi_rdata_24,afi_rdata_23,afi_rdata_22,afi_rdata_21,afi_rdata_20,afi_rdata_19,afi_rdata_18,afi_rdata_17,
afi_rdata_16,afi_rdata_15,afi_rdata_14,afi_rdata_13,afi_rdata_12,afi_rdata_11,afi_rdata_10,afi_rdata_9,afi_rdata_8,afi_rdata_7,afi_rdata_6,afi_rdata_5,afi_rdata_4,afi_rdata_3,afi_rdata_2,afi_rdata_1,afi_rdata_0}),
	.afi_wlat({afi_wlat_3,afi_wlat_2,afi_wlat_1,afi_wlat_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n({afi_cas_n_0}),
	.afi_ras_n({afi_ras_n_0}),
	.afi_rst_n({afi_rst_n_0}),
	.afi_we_n({afi_we_n_0}),
	.afi_addr({afi_addr_19,afi_addr_18,afi_addr_17,afi_addr_16,afi_addr_15,afi_addr_14,afi_addr_13,afi_addr_12,afi_addr_11,afi_addr_10,afi_addr_9,afi_addr_8,afi_addr_7,afi_addr_6,afi_addr_5,afi_addr_4,afi_addr_3,afi_addr_2,afi_addr_1,afi_addr_0}),
	.afi_ba({afi_ba_2,afi_ba_1,afi_ba_0}),
	.afi_cke({afi_cke_1,afi_cke_0}),
	.afi_cs_n({afi_cs_n_1,afi_cs_n_0}),
	.afi_dm({afi_dm_int_9,afi_dm_int_8,afi_dm_int_7,afi_dm_int_6,afi_dm_int_5,afi_dm_int_4,afi_dm_int_3,afi_dm_int_2,afi_dm_int_1,afi_dm_int_0}),
	.afi_dqs_burst({afi_dqs_burst_4,afi_dqs_burst_3,afi_dqs_burst_2,afi_dqs_burst_1,afi_dqs_burst_0}),
	.afi_odt({afi_odt_1,afi_odt_0}),
	.afi_rdata_en({afi_rdata_en_4,afi_rdata_en_3,afi_rdata_en_2,afi_rdata_en_1,afi_rdata_en_0}),
	.afi_rdata_en_full({afi_rdata_en_full_4,afi_rdata_en_full_3,afi_rdata_en_full_2,afi_rdata_en_full_1,afi_rdata_en_full_0}),
	.afi_wdata({afi_wdata_int_79,afi_wdata_int_78,afi_wdata_int_77,afi_wdata_int_76,afi_wdata_int_75,afi_wdata_int_74,afi_wdata_int_73,afi_wdata_int_72,afi_wdata_int_71,afi_wdata_int_70,afi_wdata_int_69,afi_wdata_int_68,afi_wdata_int_67,afi_wdata_int_66,afi_wdata_int_65,afi_wdata_int_64,
afi_wdata_int_63,afi_wdata_int_62,afi_wdata_int_61,afi_wdata_int_60,afi_wdata_int_59,afi_wdata_int_58,afi_wdata_int_57,afi_wdata_int_56,afi_wdata_int_55,afi_wdata_int_54,afi_wdata_int_53,afi_wdata_int_52,afi_wdata_int_51,afi_wdata_int_50,afi_wdata_int_49,afi_wdata_int_48,
afi_wdata_int_47,afi_wdata_int_46,afi_wdata_int_45,afi_wdata_int_44,afi_wdata_int_43,afi_wdata_int_42,afi_wdata_int_41,afi_wdata_int_40,afi_wdata_int_39,afi_wdata_int_38,afi_wdata_int_37,afi_wdata_int_36,afi_wdata_int_35,afi_wdata_int_34,afi_wdata_int_33,afi_wdata_int_32,
afi_wdata_int_31,afi_wdata_int_30,afi_wdata_int_29,afi_wdata_int_28,afi_wdata_int_27,afi_wdata_int_26,afi_wdata_int_25,afi_wdata_int_24,afi_wdata_int_23,afi_wdata_int_22,afi_wdata_int_21,afi_wdata_int_20,afi_wdata_int_19,afi_wdata_int_18,afi_wdata_int_17,afi_wdata_int_16,
afi_wdata_int_15,afi_wdata_int_14,afi_wdata_int_13,afi_wdata_int_12,afi_wdata_int_11,afi_wdata_int_10,afi_wdata_int_9,afi_wdata_int_8,afi_wdata_int_7,afi_wdata_int_6,afi_wdata_int_5,afi_wdata_int_4,afi_wdata_int_3,afi_wdata_int_2,afi_wdata_int_1,afi_wdata_int_0}),
	.afi_wdata_valid({afi_wdata_valid_4,afi_wdata_valid_3,afi_wdata_valid_2,afi_wdata_valid_1,afi_wdata_valid_0}),
	.cfg_addlat({gnd,gnd,gnd,cfg_addlat_wire_4,cfg_addlat_wire_3,cfg_addlat_wire_2,cfg_addlat_wire_1,cfg_addlat_wire_0}),
	.cfg_bankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth_wire_2,cfg_bankaddrwidth_wire_1,cfg_bankaddrwidth_wire_0}),
	.cfg_caswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat_wire_3,cfg_caswrlat_wire_2,cfg_caswrlat_wire_1,cfg_caswrlat_wire_0}),
	.cfg_coladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth_wire_4,cfg_coladdrwidth_wire_3,cfg_coladdrwidth_wire_2,cfg_coladdrwidth_wire_1,cfg_coladdrwidth_wire_0}),
	.cfg_csaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth_wire_2,cfg_csaddrwidth_wire_1,cfg_csaddrwidth_wire_0}),
	.cfg_devicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth_wire_3,cfg_devicewidth_wire_2,cfg_devicewidth_wire_1,cfg_devicewidth_wire_0}),
	.cfg_interfacewidth({cfg_interfacewidth_wire_7,cfg_interfacewidth_wire_6,cfg_interfacewidth_wire_5,cfg_interfacewidth_wire_4,cfg_interfacewidth_wire_3,cfg_interfacewidth_wire_2,cfg_interfacewidth_wire_1,cfg_interfacewidth_wire_0}),
	.cfg_rowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth_wire_4,cfg_rowaddrwidth_wire_3,cfg_rowaddrwidth_wire_2,cfg_rowaddrwidth_wire_1,cfg_rowaddrwidth_wire_0}),
	.cfg_tcl({gnd,gnd,gnd,cfg_tcl_wire_4,cfg_tcl_wire_3,cfg_tcl_wire_2,cfg_tcl_wire_1,cfg_tcl_wire_0}),
	.cfg_tmrd({gnd,gnd,gnd,gnd,cfg_tmrd_wire_3,cfg_tmrd_wire_2,cfg_tmrd_wire_1,cfg_tmrd_wire_0}),
	.cfg_trefi({gnd,gnd,gnd,cfg_trefi_wire_12,cfg_trefi_wire_11,cfg_trefi_wire_10,cfg_trefi_wire_9,cfg_trefi_wire_8,cfg_trefi_wire_7,cfg_trefi_wire_6,cfg_trefi_wire_5,cfg_trefi_wire_4,cfg_trefi_wire_3,cfg_trefi_wire_2,cfg_trefi_wire_1,cfg_trefi_wire_0}),
	.cfg_trfc({cfg_trfc_wire_7,cfg_trfc_wire_6,cfg_trfc_wire_5,cfg_trfc_wire_4,cfg_trfc_wire_3,cfg_trfc_wire_2,cfg_trfc_wire_1,cfg_trfc_wire_0}),
	.cfg_twr({gnd,gnd,gnd,gnd,cfg_twr_wire_3,cfg_twr_wire_2,cfg_twr_wire_1,cfg_twr_wire_0}),
	.afi_mem_clk_disable({afi_mem_clk_disable_0}),
	.cfg_dramconfig({gnd,gnd,gnd,cfg_dramconfig_wire_20,cfg_dramconfig_wire_19,cfg_dramconfig_wire_18,cfg_dramconfig_wire_17,cfg_dramconfig_wire_16,cfg_dramconfig_wire_15,cfg_dramconfig_wire_14,cfg_dramconfig_wire_13,cfg_dramconfig_wire_12,cfg_dramconfig_wire_11,cfg_dramconfig_wire_10,
cfg_dramconfig_wire_9,cfg_dramconfig_wire_8,cfg_dramconfig_wire_7,cfg_dramconfig_wire_6,cfg_dramconfig_wire_5,cfg_dramconfig_wire_4,cfg_dramconfig_wire_3,cfg_dramconfig_wire_2,cfg_dramconfig_wire_1,cfg_dramconfig_wire_0}),
	.ctl_clk(ctl_clk),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module Computer_System_hps_sdram_p0_acv_hard_memphy (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	[0:0] afi_rdata_valid;
output 	ctl_reset_n;
output 	[79:0] afi_rdata;
output 	[3:0] afi_wlat;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	[0:0] afi_cas_n;
input 	[0:0] afi_ras_n;
input 	[0:0] afi_rst_n;
input 	[0:0] afi_we_n;
input 	[19:0] afi_addr;
input 	[2:0] afi_ba;
input 	[1:0] afi_cke;
input 	[1:0] afi_cs_n;
input 	[9:0] afi_dm;
input 	[4:0] afi_dqs_burst;
input 	[1:0] afi_odt;
input 	[4:0] afi_rdata_en;
input 	[4:0] afi_rdata_en_full;
input 	[79:0] afi_wdata;
input 	[4:0] afi_wdata_valid;
input 	[7:0] cfg_addlat;
input 	[7:0] cfg_bankaddrwidth;
input 	[7:0] cfg_caswrlat;
input 	[7:0] cfg_coladdrwidth;
input 	[7:0] cfg_csaddrwidth;
input 	[7:0] cfg_devicewidth;
input 	[7:0] cfg_interfacewidth;
input 	[7:0] cfg_rowaddrwidth;
input 	[7:0] cfg_tcl;
input 	[7:0] cfg_tmrd;
input 	[15:0] cfg_trefi;
input 	[7:0] cfg_trfc;
input 	[7:0] cfg_twr;
input 	[0:0] afi_mem_clk_disable;
input 	[23:0] cfg_dramconfig;
output 	ctl_clk;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \memphy_ldc|leveled_hr_clocks[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \phy_ddio_address[0] ;
wire \phy_ddio_address[1] ;
wire \phy_ddio_address[2] ;
wire \phy_ddio_address[3] ;
wire \phy_ddio_address[4] ;
wire \phy_ddio_address[5] ;
wire \phy_ddio_address[6] ;
wire \phy_ddio_address[7] ;
wire \phy_ddio_address[8] ;
wire \phy_ddio_address[9] ;
wire \phy_ddio_address[10] ;
wire \phy_ddio_address[11] ;
wire \phy_ddio_address[12] ;
wire \phy_ddio_address[13] ;
wire \phy_ddio_address[14] ;
wire \phy_ddio_address[15] ;
wire \phy_ddio_address[16] ;
wire \phy_ddio_address[17] ;
wire \phy_ddio_address[18] ;
wire \phy_ddio_address[19] ;
wire \phy_ddio_address[20] ;
wire \phy_ddio_address[21] ;
wire \phy_ddio_address[22] ;
wire \phy_ddio_address[23] ;
wire \phy_ddio_address[24] ;
wire \phy_ddio_address[25] ;
wire \phy_ddio_address[26] ;
wire \phy_ddio_address[27] ;
wire \phy_ddio_address[28] ;
wire \phy_ddio_address[29] ;
wire \phy_ddio_address[30] ;
wire \phy_ddio_address[31] ;
wire \phy_ddio_address[32] ;
wire \phy_ddio_address[33] ;
wire \phy_ddio_address[34] ;
wire \phy_ddio_address[35] ;
wire \phy_ddio_address[36] ;
wire \phy_ddio_address[37] ;
wire \phy_ddio_address[38] ;
wire \phy_ddio_address[39] ;
wire \phy_ddio_address[40] ;
wire \phy_ddio_address[41] ;
wire \phy_ddio_address[42] ;
wire \phy_ddio_address[43] ;
wire \phy_ddio_address[44] ;
wire \phy_ddio_address[45] ;
wire \phy_ddio_address[46] ;
wire \phy_ddio_address[47] ;
wire \phy_ddio_address[48] ;
wire \phy_ddio_address[49] ;
wire \phy_ddio_address[50] ;
wire \phy_ddio_address[51] ;
wire \phy_ddio_address[52] ;
wire \phy_ddio_address[53] ;
wire \phy_ddio_address[54] ;
wire \phy_ddio_address[55] ;
wire \phy_ddio_address[56] ;
wire \phy_ddio_address[57] ;
wire \phy_ddio_address[58] ;
wire \phy_ddio_address[59] ;
wire \phy_ddio_bank[0] ;
wire \phy_ddio_bank[1] ;
wire \phy_ddio_bank[2] ;
wire \phy_ddio_bank[3] ;
wire \phy_ddio_bank[4] ;
wire \phy_ddio_bank[5] ;
wire \phy_ddio_bank[6] ;
wire \phy_ddio_bank[7] ;
wire \phy_ddio_bank[8] ;
wire \phy_ddio_bank[9] ;
wire \phy_ddio_bank[10] ;
wire \phy_ddio_bank[11] ;
wire \phy_ddio_cas_n[0] ;
wire \phy_ddio_cas_n[1] ;
wire \phy_ddio_cas_n[2] ;
wire \phy_ddio_cas_n[3] ;
wire \phy_ddio_ck[0] ;
wire \phy_ddio_ck[1] ;
wire \phy_ddio_cke[0] ;
wire \phy_ddio_cke[1] ;
wire \phy_ddio_cke[2] ;
wire \phy_ddio_cke[3] ;
wire \phy_ddio_cs_n[0] ;
wire \phy_ddio_cs_n[1] ;
wire \phy_ddio_cs_n[2] ;
wire \phy_ddio_cs_n[3] ;
wire \phy_ddio_dmdout[0] ;
wire \phy_ddio_dmdout[1] ;
wire \phy_ddio_dmdout[2] ;
wire \phy_ddio_dmdout[3] ;
wire \phy_ddio_dmdout[4] ;
wire \phy_ddio_dmdout[5] ;
wire \phy_ddio_dmdout[6] ;
wire \phy_ddio_dmdout[7] ;
wire \phy_ddio_dmdout[8] ;
wire \phy_ddio_dmdout[9] ;
wire \phy_ddio_dmdout[10] ;
wire \phy_ddio_dmdout[11] ;
wire \phy_ddio_dmdout[12] ;
wire \phy_ddio_dmdout[13] ;
wire \phy_ddio_dmdout[14] ;
wire \phy_ddio_dmdout[15] ;
wire \phy_ddio_dqdout[0] ;
wire \phy_ddio_dqdout[1] ;
wire \phy_ddio_dqdout[2] ;
wire \phy_ddio_dqdout[3] ;
wire \phy_ddio_dqdout[4] ;
wire \phy_ddio_dqdout[5] ;
wire \phy_ddio_dqdout[6] ;
wire \phy_ddio_dqdout[7] ;
wire \phy_ddio_dqdout[8] ;
wire \phy_ddio_dqdout[9] ;
wire \phy_ddio_dqdout[10] ;
wire \phy_ddio_dqdout[11] ;
wire \phy_ddio_dqdout[12] ;
wire \phy_ddio_dqdout[13] ;
wire \phy_ddio_dqdout[14] ;
wire \phy_ddio_dqdout[15] ;
wire \phy_ddio_dqdout[16] ;
wire \phy_ddio_dqdout[17] ;
wire \phy_ddio_dqdout[18] ;
wire \phy_ddio_dqdout[19] ;
wire \phy_ddio_dqdout[20] ;
wire \phy_ddio_dqdout[21] ;
wire \phy_ddio_dqdout[22] ;
wire \phy_ddio_dqdout[23] ;
wire \phy_ddio_dqdout[24] ;
wire \phy_ddio_dqdout[25] ;
wire \phy_ddio_dqdout[26] ;
wire \phy_ddio_dqdout[27] ;
wire \phy_ddio_dqdout[28] ;
wire \phy_ddio_dqdout[29] ;
wire \phy_ddio_dqdout[30] ;
wire \phy_ddio_dqdout[31] ;
wire \phy_ddio_dqdout[36] ;
wire \phy_ddio_dqdout[37] ;
wire \phy_ddio_dqdout[38] ;
wire \phy_ddio_dqdout[39] ;
wire \phy_ddio_dqdout[40] ;
wire \phy_ddio_dqdout[41] ;
wire \phy_ddio_dqdout[42] ;
wire \phy_ddio_dqdout[43] ;
wire \phy_ddio_dqdout[44] ;
wire \phy_ddio_dqdout[45] ;
wire \phy_ddio_dqdout[46] ;
wire \phy_ddio_dqdout[47] ;
wire \phy_ddio_dqdout[48] ;
wire \phy_ddio_dqdout[49] ;
wire \phy_ddio_dqdout[50] ;
wire \phy_ddio_dqdout[51] ;
wire \phy_ddio_dqdout[52] ;
wire \phy_ddio_dqdout[53] ;
wire \phy_ddio_dqdout[54] ;
wire \phy_ddio_dqdout[55] ;
wire \phy_ddio_dqdout[56] ;
wire \phy_ddio_dqdout[57] ;
wire \phy_ddio_dqdout[58] ;
wire \phy_ddio_dqdout[59] ;
wire \phy_ddio_dqdout[60] ;
wire \phy_ddio_dqdout[61] ;
wire \phy_ddio_dqdout[62] ;
wire \phy_ddio_dqdout[63] ;
wire \phy_ddio_dqdout[64] ;
wire \phy_ddio_dqdout[65] ;
wire \phy_ddio_dqdout[66] ;
wire \phy_ddio_dqdout[67] ;
wire \phy_ddio_dqdout[72] ;
wire \phy_ddio_dqdout[73] ;
wire \phy_ddio_dqdout[74] ;
wire \phy_ddio_dqdout[75] ;
wire \phy_ddio_dqdout[76] ;
wire \phy_ddio_dqdout[77] ;
wire \phy_ddio_dqdout[78] ;
wire \phy_ddio_dqdout[79] ;
wire \phy_ddio_dqdout[80] ;
wire \phy_ddio_dqdout[81] ;
wire \phy_ddio_dqdout[82] ;
wire \phy_ddio_dqdout[83] ;
wire \phy_ddio_dqdout[84] ;
wire \phy_ddio_dqdout[85] ;
wire \phy_ddio_dqdout[86] ;
wire \phy_ddio_dqdout[87] ;
wire \phy_ddio_dqdout[88] ;
wire \phy_ddio_dqdout[89] ;
wire \phy_ddio_dqdout[90] ;
wire \phy_ddio_dqdout[91] ;
wire \phy_ddio_dqdout[92] ;
wire \phy_ddio_dqdout[93] ;
wire \phy_ddio_dqdout[94] ;
wire \phy_ddio_dqdout[95] ;
wire \phy_ddio_dqdout[96] ;
wire \phy_ddio_dqdout[97] ;
wire \phy_ddio_dqdout[98] ;
wire \phy_ddio_dqdout[99] ;
wire \phy_ddio_dqdout[100] ;
wire \phy_ddio_dqdout[101] ;
wire \phy_ddio_dqdout[102] ;
wire \phy_ddio_dqdout[103] ;
wire \phy_ddio_dqdout[108] ;
wire \phy_ddio_dqdout[109] ;
wire \phy_ddio_dqdout[110] ;
wire \phy_ddio_dqdout[111] ;
wire \phy_ddio_dqdout[112] ;
wire \phy_ddio_dqdout[113] ;
wire \phy_ddio_dqdout[114] ;
wire \phy_ddio_dqdout[115] ;
wire \phy_ddio_dqdout[116] ;
wire \phy_ddio_dqdout[117] ;
wire \phy_ddio_dqdout[118] ;
wire \phy_ddio_dqdout[119] ;
wire \phy_ddio_dqdout[120] ;
wire \phy_ddio_dqdout[121] ;
wire \phy_ddio_dqdout[122] ;
wire \phy_ddio_dqdout[123] ;
wire \phy_ddio_dqdout[124] ;
wire \phy_ddio_dqdout[125] ;
wire \phy_ddio_dqdout[126] ;
wire \phy_ddio_dqdout[127] ;
wire \phy_ddio_dqdout[128] ;
wire \phy_ddio_dqdout[129] ;
wire \phy_ddio_dqdout[130] ;
wire \phy_ddio_dqdout[131] ;
wire \phy_ddio_dqdout[132] ;
wire \phy_ddio_dqdout[133] ;
wire \phy_ddio_dqdout[134] ;
wire \phy_ddio_dqdout[135] ;
wire \phy_ddio_dqdout[136] ;
wire \phy_ddio_dqdout[137] ;
wire \phy_ddio_dqdout[138] ;
wire \phy_ddio_dqdout[139] ;
wire \phy_ddio_dqoe[0] ;
wire \phy_ddio_dqoe[1] ;
wire \phy_ddio_dqoe[2] ;
wire \phy_ddio_dqoe[3] ;
wire \phy_ddio_dqoe[4] ;
wire \phy_ddio_dqoe[5] ;
wire \phy_ddio_dqoe[6] ;
wire \phy_ddio_dqoe[7] ;
wire \phy_ddio_dqoe[8] ;
wire \phy_ddio_dqoe[9] ;
wire \phy_ddio_dqoe[10] ;
wire \phy_ddio_dqoe[11] ;
wire \phy_ddio_dqoe[12] ;
wire \phy_ddio_dqoe[13] ;
wire \phy_ddio_dqoe[14] ;
wire \phy_ddio_dqoe[15] ;
wire \phy_ddio_dqoe[18] ;
wire \phy_ddio_dqoe[19] ;
wire \phy_ddio_dqoe[20] ;
wire \phy_ddio_dqoe[21] ;
wire \phy_ddio_dqoe[22] ;
wire \phy_ddio_dqoe[23] ;
wire \phy_ddio_dqoe[24] ;
wire \phy_ddio_dqoe[25] ;
wire \phy_ddio_dqoe[26] ;
wire \phy_ddio_dqoe[27] ;
wire \phy_ddio_dqoe[28] ;
wire \phy_ddio_dqoe[29] ;
wire \phy_ddio_dqoe[30] ;
wire \phy_ddio_dqoe[31] ;
wire \phy_ddio_dqoe[32] ;
wire \phy_ddio_dqoe[33] ;
wire \phy_ddio_dqoe[36] ;
wire \phy_ddio_dqoe[37] ;
wire \phy_ddio_dqoe[38] ;
wire \phy_ddio_dqoe[39] ;
wire \phy_ddio_dqoe[40] ;
wire \phy_ddio_dqoe[41] ;
wire \phy_ddio_dqoe[42] ;
wire \phy_ddio_dqoe[43] ;
wire \phy_ddio_dqoe[44] ;
wire \phy_ddio_dqoe[45] ;
wire \phy_ddio_dqoe[46] ;
wire \phy_ddio_dqoe[47] ;
wire \phy_ddio_dqoe[48] ;
wire \phy_ddio_dqoe[49] ;
wire \phy_ddio_dqoe[50] ;
wire \phy_ddio_dqoe[51] ;
wire \phy_ddio_dqoe[54] ;
wire \phy_ddio_dqoe[55] ;
wire \phy_ddio_dqoe[56] ;
wire \phy_ddio_dqoe[57] ;
wire \phy_ddio_dqoe[58] ;
wire \phy_ddio_dqoe[59] ;
wire \phy_ddio_dqoe[60] ;
wire \phy_ddio_dqoe[61] ;
wire \phy_ddio_dqoe[62] ;
wire \phy_ddio_dqoe[63] ;
wire \phy_ddio_dqoe[64] ;
wire \phy_ddio_dqoe[65] ;
wire \phy_ddio_dqoe[66] ;
wire \phy_ddio_dqoe[67] ;
wire \phy_ddio_dqoe[68] ;
wire \phy_ddio_dqoe[69] ;
wire \phy_ddio_dqs_dout[0] ;
wire \phy_ddio_dqs_dout[1] ;
wire \phy_ddio_dqs_dout[2] ;
wire \phy_ddio_dqs_dout[3] ;
wire \phy_ddio_dqs_dout[4] ;
wire \phy_ddio_dqs_dout[5] ;
wire \phy_ddio_dqs_dout[6] ;
wire \phy_ddio_dqs_dout[7] ;
wire \phy_ddio_dqs_dout[8] ;
wire \phy_ddio_dqs_dout[9] ;
wire \phy_ddio_dqs_dout[10] ;
wire \phy_ddio_dqs_dout[11] ;
wire \phy_ddio_dqs_dout[12] ;
wire \phy_ddio_dqs_dout[13] ;
wire \phy_ddio_dqs_dout[14] ;
wire \phy_ddio_dqs_dout[15] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[0] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[1] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[2] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[3] ;
wire \phy_ddio_dqslogic_aclr_pstamble[0] ;
wire \phy_ddio_dqslogic_aclr_pstamble[1] ;
wire \phy_ddio_dqslogic_aclr_pstamble[2] ;
wire \phy_ddio_dqslogic_aclr_pstamble[3] ;
wire \phy_ddio_dqslogic_dqsena[0] ;
wire \phy_ddio_dqslogic_dqsena[1] ;
wire \phy_ddio_dqslogic_dqsena[2] ;
wire \phy_ddio_dqslogic_dqsena[3] ;
wire \phy_ddio_dqslogic_dqsena[4] ;
wire \phy_ddio_dqslogic_dqsena[5] ;
wire \phy_ddio_dqslogic_dqsena[6] ;
wire \phy_ddio_dqslogic_dqsena[7] ;
wire \phy_ddio_dqslogic_fiforeset[0] ;
wire \phy_ddio_dqslogic_fiforeset[1] ;
wire \phy_ddio_dqslogic_fiforeset[2] ;
wire \phy_ddio_dqslogic_fiforeset[3] ;
wire \phy_ddio_dqslogic_incrdataen[0] ;
wire \phy_ddio_dqslogic_incrdataen[1] ;
wire \phy_ddio_dqslogic_incrdataen[2] ;
wire \phy_ddio_dqslogic_incrdataen[3] ;
wire \phy_ddio_dqslogic_incrdataen[4] ;
wire \phy_ddio_dqslogic_incrdataen[5] ;
wire \phy_ddio_dqslogic_incrdataen[6] ;
wire \phy_ddio_dqslogic_incrdataen[7] ;
wire \phy_ddio_dqslogic_incwrptr[0] ;
wire \phy_ddio_dqslogic_incwrptr[1] ;
wire \phy_ddio_dqslogic_incwrptr[2] ;
wire \phy_ddio_dqslogic_incwrptr[3] ;
wire \phy_ddio_dqslogic_incwrptr[4] ;
wire \phy_ddio_dqslogic_incwrptr[5] ;
wire \phy_ddio_dqslogic_incwrptr[6] ;
wire \phy_ddio_dqslogic_incwrptr[7] ;
wire \phy_ddio_dqslogic_oct[0] ;
wire \phy_ddio_dqslogic_oct[1] ;
wire \phy_ddio_dqslogic_oct[2] ;
wire \phy_ddio_dqslogic_oct[3] ;
wire \phy_ddio_dqslogic_oct[4] ;
wire \phy_ddio_dqslogic_oct[5] ;
wire \phy_ddio_dqslogic_oct[6] ;
wire \phy_ddio_dqslogic_oct[7] ;
wire \phy_ddio_dqslogic_readlatency[0] ;
wire \phy_ddio_dqslogic_readlatency[1] ;
wire \phy_ddio_dqslogic_readlatency[2] ;
wire \phy_ddio_dqslogic_readlatency[3] ;
wire \phy_ddio_dqslogic_readlatency[4] ;
wire \phy_ddio_dqslogic_readlatency[5] ;
wire \phy_ddio_dqslogic_readlatency[6] ;
wire \phy_ddio_dqslogic_readlatency[7] ;
wire \phy_ddio_dqslogic_readlatency[8] ;
wire \phy_ddio_dqslogic_readlatency[9] ;
wire \phy_ddio_dqslogic_readlatency[10] ;
wire \phy_ddio_dqslogic_readlatency[11] ;
wire \phy_ddio_dqslogic_readlatency[12] ;
wire \phy_ddio_dqslogic_readlatency[13] ;
wire \phy_ddio_dqslogic_readlatency[14] ;
wire \phy_ddio_dqslogic_readlatency[15] ;
wire \phy_ddio_dqslogic_readlatency[16] ;
wire \phy_ddio_dqslogic_readlatency[17] ;
wire \phy_ddio_dqslogic_readlatency[18] ;
wire \phy_ddio_dqslogic_readlatency[19] ;
wire \phy_ddio_dqs_oe[0] ;
wire \phy_ddio_dqs_oe[1] ;
wire \phy_ddio_dqs_oe[2] ;
wire \phy_ddio_dqs_oe[3] ;
wire \phy_ddio_dqs_oe[4] ;
wire \phy_ddio_dqs_oe[5] ;
wire \phy_ddio_dqs_oe[6] ;
wire \phy_ddio_dqs_oe[7] ;
wire \phy_ddio_odt[0] ;
wire \phy_ddio_odt[1] ;
wire \phy_ddio_odt[2] ;
wire \phy_ddio_odt[3] ;
wire \phy_ddio_ras_n[0] ;
wire \phy_ddio_ras_n[1] ;
wire \phy_ddio_ras_n[2] ;
wire \phy_ddio_ras_n[3] ;
wire \phy_ddio_reset_n[0] ;
wire \phy_ddio_reset_n[1] ;
wire \phy_ddio_reset_n[2] ;
wire \phy_ddio_reset_n[3] ;
wire \phy_ddio_we_n[0] ;
wire \phy_ddio_we_n[1] ;
wire \phy_ddio_we_n[2] ;
wire \phy_ddio_we_n[3] ;

wire [79:0] hphy_inst_AFIRDATA_bus;
wire [3:0] hphy_inst_AFIWLAT_bus;
wire [63:0] hphy_inst_PHYDDIOADDRDOUT_bus;
wire [11:0] hphy_inst_PHYDDIOBADOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCKDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCKEDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCSNDOUT_bus;
wire [19:0] hphy_inst_PHYDDIODMDOUT_bus;
wire [179:0] hphy_inst_PHYDDIODQDOUT_bus;
wire [89:0] hphy_inst_PHYDDIODQOE_bus;
wire [19:0] hphy_inst_PHYDDIODQSDOUT_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICDQSENA_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICFIFORESET_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICOCT_bus;
wire [24:0] hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus;
wire [9:0] hphy_inst_PHYDDIODQSOE_bus;
wire [7:0] hphy_inst_PHYDDIOODTDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORESETNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOWENDOUT_bus;

assign afi_rdata[0] = hphy_inst_AFIRDATA_bus[0];
assign afi_rdata[1] = hphy_inst_AFIRDATA_bus[1];
assign afi_rdata[2] = hphy_inst_AFIRDATA_bus[2];
assign afi_rdata[3] = hphy_inst_AFIRDATA_bus[3];
assign afi_rdata[4] = hphy_inst_AFIRDATA_bus[4];
assign afi_rdata[5] = hphy_inst_AFIRDATA_bus[5];
assign afi_rdata[6] = hphy_inst_AFIRDATA_bus[6];
assign afi_rdata[7] = hphy_inst_AFIRDATA_bus[7];
assign afi_rdata[8] = hphy_inst_AFIRDATA_bus[8];
assign afi_rdata[9] = hphy_inst_AFIRDATA_bus[9];
assign afi_rdata[10] = hphy_inst_AFIRDATA_bus[10];
assign afi_rdata[11] = hphy_inst_AFIRDATA_bus[11];
assign afi_rdata[12] = hphy_inst_AFIRDATA_bus[12];
assign afi_rdata[13] = hphy_inst_AFIRDATA_bus[13];
assign afi_rdata[14] = hphy_inst_AFIRDATA_bus[14];
assign afi_rdata[15] = hphy_inst_AFIRDATA_bus[15];
assign afi_rdata[16] = hphy_inst_AFIRDATA_bus[16];
assign afi_rdata[17] = hphy_inst_AFIRDATA_bus[17];
assign afi_rdata[18] = hphy_inst_AFIRDATA_bus[18];
assign afi_rdata[19] = hphy_inst_AFIRDATA_bus[19];
assign afi_rdata[20] = hphy_inst_AFIRDATA_bus[20];
assign afi_rdata[21] = hphy_inst_AFIRDATA_bus[21];
assign afi_rdata[22] = hphy_inst_AFIRDATA_bus[22];
assign afi_rdata[23] = hphy_inst_AFIRDATA_bus[23];
assign afi_rdata[24] = hphy_inst_AFIRDATA_bus[24];
assign afi_rdata[25] = hphy_inst_AFIRDATA_bus[25];
assign afi_rdata[26] = hphy_inst_AFIRDATA_bus[26];
assign afi_rdata[27] = hphy_inst_AFIRDATA_bus[27];
assign afi_rdata[28] = hphy_inst_AFIRDATA_bus[28];
assign afi_rdata[29] = hphy_inst_AFIRDATA_bus[29];
assign afi_rdata[30] = hphy_inst_AFIRDATA_bus[30];
assign afi_rdata[31] = hphy_inst_AFIRDATA_bus[31];
assign afi_rdata[32] = hphy_inst_AFIRDATA_bus[32];
assign afi_rdata[33] = hphy_inst_AFIRDATA_bus[33];
assign afi_rdata[34] = hphy_inst_AFIRDATA_bus[34];
assign afi_rdata[35] = hphy_inst_AFIRDATA_bus[35];
assign afi_rdata[36] = hphy_inst_AFIRDATA_bus[36];
assign afi_rdata[37] = hphy_inst_AFIRDATA_bus[37];
assign afi_rdata[38] = hphy_inst_AFIRDATA_bus[38];
assign afi_rdata[39] = hphy_inst_AFIRDATA_bus[39];
assign afi_rdata[40] = hphy_inst_AFIRDATA_bus[40];
assign afi_rdata[41] = hphy_inst_AFIRDATA_bus[41];
assign afi_rdata[42] = hphy_inst_AFIRDATA_bus[42];
assign afi_rdata[43] = hphy_inst_AFIRDATA_bus[43];
assign afi_rdata[44] = hphy_inst_AFIRDATA_bus[44];
assign afi_rdata[45] = hphy_inst_AFIRDATA_bus[45];
assign afi_rdata[46] = hphy_inst_AFIRDATA_bus[46];
assign afi_rdata[47] = hphy_inst_AFIRDATA_bus[47];
assign afi_rdata[48] = hphy_inst_AFIRDATA_bus[48];
assign afi_rdata[49] = hphy_inst_AFIRDATA_bus[49];
assign afi_rdata[50] = hphy_inst_AFIRDATA_bus[50];
assign afi_rdata[51] = hphy_inst_AFIRDATA_bus[51];
assign afi_rdata[52] = hphy_inst_AFIRDATA_bus[52];
assign afi_rdata[53] = hphy_inst_AFIRDATA_bus[53];
assign afi_rdata[54] = hphy_inst_AFIRDATA_bus[54];
assign afi_rdata[55] = hphy_inst_AFIRDATA_bus[55];
assign afi_rdata[56] = hphy_inst_AFIRDATA_bus[56];
assign afi_rdata[57] = hphy_inst_AFIRDATA_bus[57];
assign afi_rdata[58] = hphy_inst_AFIRDATA_bus[58];
assign afi_rdata[59] = hphy_inst_AFIRDATA_bus[59];
assign afi_rdata[60] = hphy_inst_AFIRDATA_bus[60];
assign afi_rdata[61] = hphy_inst_AFIRDATA_bus[61];
assign afi_rdata[62] = hphy_inst_AFIRDATA_bus[62];
assign afi_rdata[63] = hphy_inst_AFIRDATA_bus[63];
assign afi_rdata[64] = hphy_inst_AFIRDATA_bus[64];
assign afi_rdata[65] = hphy_inst_AFIRDATA_bus[65];
assign afi_rdata[66] = hphy_inst_AFIRDATA_bus[66];
assign afi_rdata[67] = hphy_inst_AFIRDATA_bus[67];
assign afi_rdata[68] = hphy_inst_AFIRDATA_bus[68];
assign afi_rdata[69] = hphy_inst_AFIRDATA_bus[69];
assign afi_rdata[70] = hphy_inst_AFIRDATA_bus[70];
assign afi_rdata[71] = hphy_inst_AFIRDATA_bus[71];
assign afi_rdata[72] = hphy_inst_AFIRDATA_bus[72];
assign afi_rdata[73] = hphy_inst_AFIRDATA_bus[73];
assign afi_rdata[74] = hphy_inst_AFIRDATA_bus[74];
assign afi_rdata[75] = hphy_inst_AFIRDATA_bus[75];
assign afi_rdata[76] = hphy_inst_AFIRDATA_bus[76];
assign afi_rdata[77] = hphy_inst_AFIRDATA_bus[77];
assign afi_rdata[78] = hphy_inst_AFIRDATA_bus[78];
assign afi_rdata[79] = hphy_inst_AFIRDATA_bus[79];

assign afi_wlat[0] = hphy_inst_AFIWLAT_bus[0];
assign afi_wlat[1] = hphy_inst_AFIWLAT_bus[1];
assign afi_wlat[2] = hphy_inst_AFIWLAT_bus[2];
assign afi_wlat[3] = hphy_inst_AFIWLAT_bus[3];

assign \phy_ddio_address[0]  = hphy_inst_PHYDDIOADDRDOUT_bus[0];
assign \phy_ddio_address[1]  = hphy_inst_PHYDDIOADDRDOUT_bus[1];
assign \phy_ddio_address[2]  = hphy_inst_PHYDDIOADDRDOUT_bus[2];
assign \phy_ddio_address[3]  = hphy_inst_PHYDDIOADDRDOUT_bus[3];
assign \phy_ddio_address[4]  = hphy_inst_PHYDDIOADDRDOUT_bus[4];
assign \phy_ddio_address[5]  = hphy_inst_PHYDDIOADDRDOUT_bus[5];
assign \phy_ddio_address[6]  = hphy_inst_PHYDDIOADDRDOUT_bus[6];
assign \phy_ddio_address[7]  = hphy_inst_PHYDDIOADDRDOUT_bus[7];
assign \phy_ddio_address[8]  = hphy_inst_PHYDDIOADDRDOUT_bus[8];
assign \phy_ddio_address[9]  = hphy_inst_PHYDDIOADDRDOUT_bus[9];
assign \phy_ddio_address[10]  = hphy_inst_PHYDDIOADDRDOUT_bus[10];
assign \phy_ddio_address[11]  = hphy_inst_PHYDDIOADDRDOUT_bus[11];
assign \phy_ddio_address[12]  = hphy_inst_PHYDDIOADDRDOUT_bus[12];
assign \phy_ddio_address[13]  = hphy_inst_PHYDDIOADDRDOUT_bus[13];
assign \phy_ddio_address[14]  = hphy_inst_PHYDDIOADDRDOUT_bus[14];
assign \phy_ddio_address[15]  = hphy_inst_PHYDDIOADDRDOUT_bus[15];
assign \phy_ddio_address[16]  = hphy_inst_PHYDDIOADDRDOUT_bus[16];
assign \phy_ddio_address[17]  = hphy_inst_PHYDDIOADDRDOUT_bus[17];
assign \phy_ddio_address[18]  = hphy_inst_PHYDDIOADDRDOUT_bus[18];
assign \phy_ddio_address[19]  = hphy_inst_PHYDDIOADDRDOUT_bus[19];
assign \phy_ddio_address[20]  = hphy_inst_PHYDDIOADDRDOUT_bus[20];
assign \phy_ddio_address[21]  = hphy_inst_PHYDDIOADDRDOUT_bus[21];
assign \phy_ddio_address[22]  = hphy_inst_PHYDDIOADDRDOUT_bus[22];
assign \phy_ddio_address[23]  = hphy_inst_PHYDDIOADDRDOUT_bus[23];
assign \phy_ddio_address[24]  = hphy_inst_PHYDDIOADDRDOUT_bus[24];
assign \phy_ddio_address[25]  = hphy_inst_PHYDDIOADDRDOUT_bus[25];
assign \phy_ddio_address[26]  = hphy_inst_PHYDDIOADDRDOUT_bus[26];
assign \phy_ddio_address[27]  = hphy_inst_PHYDDIOADDRDOUT_bus[27];
assign \phy_ddio_address[28]  = hphy_inst_PHYDDIOADDRDOUT_bus[28];
assign \phy_ddio_address[29]  = hphy_inst_PHYDDIOADDRDOUT_bus[29];
assign \phy_ddio_address[30]  = hphy_inst_PHYDDIOADDRDOUT_bus[30];
assign \phy_ddio_address[31]  = hphy_inst_PHYDDIOADDRDOUT_bus[31];
assign \phy_ddio_address[32]  = hphy_inst_PHYDDIOADDRDOUT_bus[32];
assign \phy_ddio_address[33]  = hphy_inst_PHYDDIOADDRDOUT_bus[33];
assign \phy_ddio_address[34]  = hphy_inst_PHYDDIOADDRDOUT_bus[34];
assign \phy_ddio_address[35]  = hphy_inst_PHYDDIOADDRDOUT_bus[35];
assign \phy_ddio_address[36]  = hphy_inst_PHYDDIOADDRDOUT_bus[36];
assign \phy_ddio_address[37]  = hphy_inst_PHYDDIOADDRDOUT_bus[37];
assign \phy_ddio_address[38]  = hphy_inst_PHYDDIOADDRDOUT_bus[38];
assign \phy_ddio_address[39]  = hphy_inst_PHYDDIOADDRDOUT_bus[39];
assign \phy_ddio_address[40]  = hphy_inst_PHYDDIOADDRDOUT_bus[40];
assign \phy_ddio_address[41]  = hphy_inst_PHYDDIOADDRDOUT_bus[41];
assign \phy_ddio_address[42]  = hphy_inst_PHYDDIOADDRDOUT_bus[42];
assign \phy_ddio_address[43]  = hphy_inst_PHYDDIOADDRDOUT_bus[43];
assign \phy_ddio_address[44]  = hphy_inst_PHYDDIOADDRDOUT_bus[44];
assign \phy_ddio_address[45]  = hphy_inst_PHYDDIOADDRDOUT_bus[45];
assign \phy_ddio_address[46]  = hphy_inst_PHYDDIOADDRDOUT_bus[46];
assign \phy_ddio_address[47]  = hphy_inst_PHYDDIOADDRDOUT_bus[47];
assign \phy_ddio_address[48]  = hphy_inst_PHYDDIOADDRDOUT_bus[48];
assign \phy_ddio_address[49]  = hphy_inst_PHYDDIOADDRDOUT_bus[49];
assign \phy_ddio_address[50]  = hphy_inst_PHYDDIOADDRDOUT_bus[50];
assign \phy_ddio_address[51]  = hphy_inst_PHYDDIOADDRDOUT_bus[51];
assign \phy_ddio_address[52]  = hphy_inst_PHYDDIOADDRDOUT_bus[52];
assign \phy_ddio_address[53]  = hphy_inst_PHYDDIOADDRDOUT_bus[53];
assign \phy_ddio_address[54]  = hphy_inst_PHYDDIOADDRDOUT_bus[54];
assign \phy_ddio_address[55]  = hphy_inst_PHYDDIOADDRDOUT_bus[55];
assign \phy_ddio_address[56]  = hphy_inst_PHYDDIOADDRDOUT_bus[56];
assign \phy_ddio_address[57]  = hphy_inst_PHYDDIOADDRDOUT_bus[57];
assign \phy_ddio_address[58]  = hphy_inst_PHYDDIOADDRDOUT_bus[58];
assign \phy_ddio_address[59]  = hphy_inst_PHYDDIOADDRDOUT_bus[59];

assign \phy_ddio_bank[0]  = hphy_inst_PHYDDIOBADOUT_bus[0];
assign \phy_ddio_bank[1]  = hphy_inst_PHYDDIOBADOUT_bus[1];
assign \phy_ddio_bank[2]  = hphy_inst_PHYDDIOBADOUT_bus[2];
assign \phy_ddio_bank[3]  = hphy_inst_PHYDDIOBADOUT_bus[3];
assign \phy_ddio_bank[4]  = hphy_inst_PHYDDIOBADOUT_bus[4];
assign \phy_ddio_bank[5]  = hphy_inst_PHYDDIOBADOUT_bus[5];
assign \phy_ddio_bank[6]  = hphy_inst_PHYDDIOBADOUT_bus[6];
assign \phy_ddio_bank[7]  = hphy_inst_PHYDDIOBADOUT_bus[7];
assign \phy_ddio_bank[8]  = hphy_inst_PHYDDIOBADOUT_bus[8];
assign \phy_ddio_bank[9]  = hphy_inst_PHYDDIOBADOUT_bus[9];
assign \phy_ddio_bank[10]  = hphy_inst_PHYDDIOBADOUT_bus[10];
assign \phy_ddio_bank[11]  = hphy_inst_PHYDDIOBADOUT_bus[11];

assign \phy_ddio_cas_n[0]  = hphy_inst_PHYDDIOCASNDOUT_bus[0];
assign \phy_ddio_cas_n[1]  = hphy_inst_PHYDDIOCASNDOUT_bus[1];
assign \phy_ddio_cas_n[2]  = hphy_inst_PHYDDIOCASNDOUT_bus[2];
assign \phy_ddio_cas_n[3]  = hphy_inst_PHYDDIOCASNDOUT_bus[3];

assign \phy_ddio_ck[0]  = hphy_inst_PHYDDIOCKDOUT_bus[0];
assign \phy_ddio_ck[1]  = hphy_inst_PHYDDIOCKDOUT_bus[1];

assign \phy_ddio_cke[0]  = hphy_inst_PHYDDIOCKEDOUT_bus[0];
assign \phy_ddio_cke[1]  = hphy_inst_PHYDDIOCKEDOUT_bus[1];
assign \phy_ddio_cke[2]  = hphy_inst_PHYDDIOCKEDOUT_bus[2];
assign \phy_ddio_cke[3]  = hphy_inst_PHYDDIOCKEDOUT_bus[3];

assign \phy_ddio_cs_n[0]  = hphy_inst_PHYDDIOCSNDOUT_bus[0];
assign \phy_ddio_cs_n[1]  = hphy_inst_PHYDDIOCSNDOUT_bus[1];
assign \phy_ddio_cs_n[2]  = hphy_inst_PHYDDIOCSNDOUT_bus[2];
assign \phy_ddio_cs_n[3]  = hphy_inst_PHYDDIOCSNDOUT_bus[3];

assign \phy_ddio_dmdout[0]  = hphy_inst_PHYDDIODMDOUT_bus[0];
assign \phy_ddio_dmdout[1]  = hphy_inst_PHYDDIODMDOUT_bus[1];
assign \phy_ddio_dmdout[2]  = hphy_inst_PHYDDIODMDOUT_bus[2];
assign \phy_ddio_dmdout[3]  = hphy_inst_PHYDDIODMDOUT_bus[3];
assign \phy_ddio_dmdout[4]  = hphy_inst_PHYDDIODMDOUT_bus[4];
assign \phy_ddio_dmdout[5]  = hphy_inst_PHYDDIODMDOUT_bus[5];
assign \phy_ddio_dmdout[6]  = hphy_inst_PHYDDIODMDOUT_bus[6];
assign \phy_ddio_dmdout[7]  = hphy_inst_PHYDDIODMDOUT_bus[7];
assign \phy_ddio_dmdout[8]  = hphy_inst_PHYDDIODMDOUT_bus[8];
assign \phy_ddio_dmdout[9]  = hphy_inst_PHYDDIODMDOUT_bus[9];
assign \phy_ddio_dmdout[10]  = hphy_inst_PHYDDIODMDOUT_bus[10];
assign \phy_ddio_dmdout[11]  = hphy_inst_PHYDDIODMDOUT_bus[11];
assign \phy_ddio_dmdout[12]  = hphy_inst_PHYDDIODMDOUT_bus[12];
assign \phy_ddio_dmdout[13]  = hphy_inst_PHYDDIODMDOUT_bus[13];
assign \phy_ddio_dmdout[14]  = hphy_inst_PHYDDIODMDOUT_bus[14];
assign \phy_ddio_dmdout[15]  = hphy_inst_PHYDDIODMDOUT_bus[15];

assign \phy_ddio_dqdout[0]  = hphy_inst_PHYDDIODQDOUT_bus[0];
assign \phy_ddio_dqdout[1]  = hphy_inst_PHYDDIODQDOUT_bus[1];
assign \phy_ddio_dqdout[2]  = hphy_inst_PHYDDIODQDOUT_bus[2];
assign \phy_ddio_dqdout[3]  = hphy_inst_PHYDDIODQDOUT_bus[3];
assign \phy_ddio_dqdout[4]  = hphy_inst_PHYDDIODQDOUT_bus[4];
assign \phy_ddio_dqdout[5]  = hphy_inst_PHYDDIODQDOUT_bus[5];
assign \phy_ddio_dqdout[6]  = hphy_inst_PHYDDIODQDOUT_bus[6];
assign \phy_ddio_dqdout[7]  = hphy_inst_PHYDDIODQDOUT_bus[7];
assign \phy_ddio_dqdout[8]  = hphy_inst_PHYDDIODQDOUT_bus[8];
assign \phy_ddio_dqdout[9]  = hphy_inst_PHYDDIODQDOUT_bus[9];
assign \phy_ddio_dqdout[10]  = hphy_inst_PHYDDIODQDOUT_bus[10];
assign \phy_ddio_dqdout[11]  = hphy_inst_PHYDDIODQDOUT_bus[11];
assign \phy_ddio_dqdout[12]  = hphy_inst_PHYDDIODQDOUT_bus[12];
assign \phy_ddio_dqdout[13]  = hphy_inst_PHYDDIODQDOUT_bus[13];
assign \phy_ddio_dqdout[14]  = hphy_inst_PHYDDIODQDOUT_bus[14];
assign \phy_ddio_dqdout[15]  = hphy_inst_PHYDDIODQDOUT_bus[15];
assign \phy_ddio_dqdout[16]  = hphy_inst_PHYDDIODQDOUT_bus[16];
assign \phy_ddio_dqdout[17]  = hphy_inst_PHYDDIODQDOUT_bus[17];
assign \phy_ddio_dqdout[18]  = hphy_inst_PHYDDIODQDOUT_bus[18];
assign \phy_ddio_dqdout[19]  = hphy_inst_PHYDDIODQDOUT_bus[19];
assign \phy_ddio_dqdout[20]  = hphy_inst_PHYDDIODQDOUT_bus[20];
assign \phy_ddio_dqdout[21]  = hphy_inst_PHYDDIODQDOUT_bus[21];
assign \phy_ddio_dqdout[22]  = hphy_inst_PHYDDIODQDOUT_bus[22];
assign \phy_ddio_dqdout[23]  = hphy_inst_PHYDDIODQDOUT_bus[23];
assign \phy_ddio_dqdout[24]  = hphy_inst_PHYDDIODQDOUT_bus[24];
assign \phy_ddio_dqdout[25]  = hphy_inst_PHYDDIODQDOUT_bus[25];
assign \phy_ddio_dqdout[26]  = hphy_inst_PHYDDIODQDOUT_bus[26];
assign \phy_ddio_dqdout[27]  = hphy_inst_PHYDDIODQDOUT_bus[27];
assign \phy_ddio_dqdout[28]  = hphy_inst_PHYDDIODQDOUT_bus[28];
assign \phy_ddio_dqdout[29]  = hphy_inst_PHYDDIODQDOUT_bus[29];
assign \phy_ddio_dqdout[30]  = hphy_inst_PHYDDIODQDOUT_bus[30];
assign \phy_ddio_dqdout[31]  = hphy_inst_PHYDDIODQDOUT_bus[31];
assign \phy_ddio_dqdout[36]  = hphy_inst_PHYDDIODQDOUT_bus[36];
assign \phy_ddio_dqdout[37]  = hphy_inst_PHYDDIODQDOUT_bus[37];
assign \phy_ddio_dqdout[38]  = hphy_inst_PHYDDIODQDOUT_bus[38];
assign \phy_ddio_dqdout[39]  = hphy_inst_PHYDDIODQDOUT_bus[39];
assign \phy_ddio_dqdout[40]  = hphy_inst_PHYDDIODQDOUT_bus[40];
assign \phy_ddio_dqdout[41]  = hphy_inst_PHYDDIODQDOUT_bus[41];
assign \phy_ddio_dqdout[42]  = hphy_inst_PHYDDIODQDOUT_bus[42];
assign \phy_ddio_dqdout[43]  = hphy_inst_PHYDDIODQDOUT_bus[43];
assign \phy_ddio_dqdout[44]  = hphy_inst_PHYDDIODQDOUT_bus[44];
assign \phy_ddio_dqdout[45]  = hphy_inst_PHYDDIODQDOUT_bus[45];
assign \phy_ddio_dqdout[46]  = hphy_inst_PHYDDIODQDOUT_bus[46];
assign \phy_ddio_dqdout[47]  = hphy_inst_PHYDDIODQDOUT_bus[47];
assign \phy_ddio_dqdout[48]  = hphy_inst_PHYDDIODQDOUT_bus[48];
assign \phy_ddio_dqdout[49]  = hphy_inst_PHYDDIODQDOUT_bus[49];
assign \phy_ddio_dqdout[50]  = hphy_inst_PHYDDIODQDOUT_bus[50];
assign \phy_ddio_dqdout[51]  = hphy_inst_PHYDDIODQDOUT_bus[51];
assign \phy_ddio_dqdout[52]  = hphy_inst_PHYDDIODQDOUT_bus[52];
assign \phy_ddio_dqdout[53]  = hphy_inst_PHYDDIODQDOUT_bus[53];
assign \phy_ddio_dqdout[54]  = hphy_inst_PHYDDIODQDOUT_bus[54];
assign \phy_ddio_dqdout[55]  = hphy_inst_PHYDDIODQDOUT_bus[55];
assign \phy_ddio_dqdout[56]  = hphy_inst_PHYDDIODQDOUT_bus[56];
assign \phy_ddio_dqdout[57]  = hphy_inst_PHYDDIODQDOUT_bus[57];
assign \phy_ddio_dqdout[58]  = hphy_inst_PHYDDIODQDOUT_bus[58];
assign \phy_ddio_dqdout[59]  = hphy_inst_PHYDDIODQDOUT_bus[59];
assign \phy_ddio_dqdout[60]  = hphy_inst_PHYDDIODQDOUT_bus[60];
assign \phy_ddio_dqdout[61]  = hphy_inst_PHYDDIODQDOUT_bus[61];
assign \phy_ddio_dqdout[62]  = hphy_inst_PHYDDIODQDOUT_bus[62];
assign \phy_ddio_dqdout[63]  = hphy_inst_PHYDDIODQDOUT_bus[63];
assign \phy_ddio_dqdout[64]  = hphy_inst_PHYDDIODQDOUT_bus[64];
assign \phy_ddio_dqdout[65]  = hphy_inst_PHYDDIODQDOUT_bus[65];
assign \phy_ddio_dqdout[66]  = hphy_inst_PHYDDIODQDOUT_bus[66];
assign \phy_ddio_dqdout[67]  = hphy_inst_PHYDDIODQDOUT_bus[67];
assign \phy_ddio_dqdout[72]  = hphy_inst_PHYDDIODQDOUT_bus[72];
assign \phy_ddio_dqdout[73]  = hphy_inst_PHYDDIODQDOUT_bus[73];
assign \phy_ddio_dqdout[74]  = hphy_inst_PHYDDIODQDOUT_bus[74];
assign \phy_ddio_dqdout[75]  = hphy_inst_PHYDDIODQDOUT_bus[75];
assign \phy_ddio_dqdout[76]  = hphy_inst_PHYDDIODQDOUT_bus[76];
assign \phy_ddio_dqdout[77]  = hphy_inst_PHYDDIODQDOUT_bus[77];
assign \phy_ddio_dqdout[78]  = hphy_inst_PHYDDIODQDOUT_bus[78];
assign \phy_ddio_dqdout[79]  = hphy_inst_PHYDDIODQDOUT_bus[79];
assign \phy_ddio_dqdout[80]  = hphy_inst_PHYDDIODQDOUT_bus[80];
assign \phy_ddio_dqdout[81]  = hphy_inst_PHYDDIODQDOUT_bus[81];
assign \phy_ddio_dqdout[82]  = hphy_inst_PHYDDIODQDOUT_bus[82];
assign \phy_ddio_dqdout[83]  = hphy_inst_PHYDDIODQDOUT_bus[83];
assign \phy_ddio_dqdout[84]  = hphy_inst_PHYDDIODQDOUT_bus[84];
assign \phy_ddio_dqdout[85]  = hphy_inst_PHYDDIODQDOUT_bus[85];
assign \phy_ddio_dqdout[86]  = hphy_inst_PHYDDIODQDOUT_bus[86];
assign \phy_ddio_dqdout[87]  = hphy_inst_PHYDDIODQDOUT_bus[87];
assign \phy_ddio_dqdout[88]  = hphy_inst_PHYDDIODQDOUT_bus[88];
assign \phy_ddio_dqdout[89]  = hphy_inst_PHYDDIODQDOUT_bus[89];
assign \phy_ddio_dqdout[90]  = hphy_inst_PHYDDIODQDOUT_bus[90];
assign \phy_ddio_dqdout[91]  = hphy_inst_PHYDDIODQDOUT_bus[91];
assign \phy_ddio_dqdout[92]  = hphy_inst_PHYDDIODQDOUT_bus[92];
assign \phy_ddio_dqdout[93]  = hphy_inst_PHYDDIODQDOUT_bus[93];
assign \phy_ddio_dqdout[94]  = hphy_inst_PHYDDIODQDOUT_bus[94];
assign \phy_ddio_dqdout[95]  = hphy_inst_PHYDDIODQDOUT_bus[95];
assign \phy_ddio_dqdout[96]  = hphy_inst_PHYDDIODQDOUT_bus[96];
assign \phy_ddio_dqdout[97]  = hphy_inst_PHYDDIODQDOUT_bus[97];
assign \phy_ddio_dqdout[98]  = hphy_inst_PHYDDIODQDOUT_bus[98];
assign \phy_ddio_dqdout[99]  = hphy_inst_PHYDDIODQDOUT_bus[99];
assign \phy_ddio_dqdout[100]  = hphy_inst_PHYDDIODQDOUT_bus[100];
assign \phy_ddio_dqdout[101]  = hphy_inst_PHYDDIODQDOUT_bus[101];
assign \phy_ddio_dqdout[102]  = hphy_inst_PHYDDIODQDOUT_bus[102];
assign \phy_ddio_dqdout[103]  = hphy_inst_PHYDDIODQDOUT_bus[103];
assign \phy_ddio_dqdout[108]  = hphy_inst_PHYDDIODQDOUT_bus[108];
assign \phy_ddio_dqdout[109]  = hphy_inst_PHYDDIODQDOUT_bus[109];
assign \phy_ddio_dqdout[110]  = hphy_inst_PHYDDIODQDOUT_bus[110];
assign \phy_ddio_dqdout[111]  = hphy_inst_PHYDDIODQDOUT_bus[111];
assign \phy_ddio_dqdout[112]  = hphy_inst_PHYDDIODQDOUT_bus[112];
assign \phy_ddio_dqdout[113]  = hphy_inst_PHYDDIODQDOUT_bus[113];
assign \phy_ddio_dqdout[114]  = hphy_inst_PHYDDIODQDOUT_bus[114];
assign \phy_ddio_dqdout[115]  = hphy_inst_PHYDDIODQDOUT_bus[115];
assign \phy_ddio_dqdout[116]  = hphy_inst_PHYDDIODQDOUT_bus[116];
assign \phy_ddio_dqdout[117]  = hphy_inst_PHYDDIODQDOUT_bus[117];
assign \phy_ddio_dqdout[118]  = hphy_inst_PHYDDIODQDOUT_bus[118];
assign \phy_ddio_dqdout[119]  = hphy_inst_PHYDDIODQDOUT_bus[119];
assign \phy_ddio_dqdout[120]  = hphy_inst_PHYDDIODQDOUT_bus[120];
assign \phy_ddio_dqdout[121]  = hphy_inst_PHYDDIODQDOUT_bus[121];
assign \phy_ddio_dqdout[122]  = hphy_inst_PHYDDIODQDOUT_bus[122];
assign \phy_ddio_dqdout[123]  = hphy_inst_PHYDDIODQDOUT_bus[123];
assign \phy_ddio_dqdout[124]  = hphy_inst_PHYDDIODQDOUT_bus[124];
assign \phy_ddio_dqdout[125]  = hphy_inst_PHYDDIODQDOUT_bus[125];
assign \phy_ddio_dqdout[126]  = hphy_inst_PHYDDIODQDOUT_bus[126];
assign \phy_ddio_dqdout[127]  = hphy_inst_PHYDDIODQDOUT_bus[127];
assign \phy_ddio_dqdout[128]  = hphy_inst_PHYDDIODQDOUT_bus[128];
assign \phy_ddio_dqdout[129]  = hphy_inst_PHYDDIODQDOUT_bus[129];
assign \phy_ddio_dqdout[130]  = hphy_inst_PHYDDIODQDOUT_bus[130];
assign \phy_ddio_dqdout[131]  = hphy_inst_PHYDDIODQDOUT_bus[131];
assign \phy_ddio_dqdout[132]  = hphy_inst_PHYDDIODQDOUT_bus[132];
assign \phy_ddio_dqdout[133]  = hphy_inst_PHYDDIODQDOUT_bus[133];
assign \phy_ddio_dqdout[134]  = hphy_inst_PHYDDIODQDOUT_bus[134];
assign \phy_ddio_dqdout[135]  = hphy_inst_PHYDDIODQDOUT_bus[135];
assign \phy_ddio_dqdout[136]  = hphy_inst_PHYDDIODQDOUT_bus[136];
assign \phy_ddio_dqdout[137]  = hphy_inst_PHYDDIODQDOUT_bus[137];
assign \phy_ddio_dqdout[138]  = hphy_inst_PHYDDIODQDOUT_bus[138];
assign \phy_ddio_dqdout[139]  = hphy_inst_PHYDDIODQDOUT_bus[139];

assign \phy_ddio_dqoe[0]  = hphy_inst_PHYDDIODQOE_bus[0];
assign \phy_ddio_dqoe[1]  = hphy_inst_PHYDDIODQOE_bus[1];
assign \phy_ddio_dqoe[2]  = hphy_inst_PHYDDIODQOE_bus[2];
assign \phy_ddio_dqoe[3]  = hphy_inst_PHYDDIODQOE_bus[3];
assign \phy_ddio_dqoe[4]  = hphy_inst_PHYDDIODQOE_bus[4];
assign \phy_ddio_dqoe[5]  = hphy_inst_PHYDDIODQOE_bus[5];
assign \phy_ddio_dqoe[6]  = hphy_inst_PHYDDIODQOE_bus[6];
assign \phy_ddio_dqoe[7]  = hphy_inst_PHYDDIODQOE_bus[7];
assign \phy_ddio_dqoe[8]  = hphy_inst_PHYDDIODQOE_bus[8];
assign \phy_ddio_dqoe[9]  = hphy_inst_PHYDDIODQOE_bus[9];
assign \phy_ddio_dqoe[10]  = hphy_inst_PHYDDIODQOE_bus[10];
assign \phy_ddio_dqoe[11]  = hphy_inst_PHYDDIODQOE_bus[11];
assign \phy_ddio_dqoe[12]  = hphy_inst_PHYDDIODQOE_bus[12];
assign \phy_ddio_dqoe[13]  = hphy_inst_PHYDDIODQOE_bus[13];
assign \phy_ddio_dqoe[14]  = hphy_inst_PHYDDIODQOE_bus[14];
assign \phy_ddio_dqoe[15]  = hphy_inst_PHYDDIODQOE_bus[15];
assign \phy_ddio_dqoe[18]  = hphy_inst_PHYDDIODQOE_bus[18];
assign \phy_ddio_dqoe[19]  = hphy_inst_PHYDDIODQOE_bus[19];
assign \phy_ddio_dqoe[20]  = hphy_inst_PHYDDIODQOE_bus[20];
assign \phy_ddio_dqoe[21]  = hphy_inst_PHYDDIODQOE_bus[21];
assign \phy_ddio_dqoe[22]  = hphy_inst_PHYDDIODQOE_bus[22];
assign \phy_ddio_dqoe[23]  = hphy_inst_PHYDDIODQOE_bus[23];
assign \phy_ddio_dqoe[24]  = hphy_inst_PHYDDIODQOE_bus[24];
assign \phy_ddio_dqoe[25]  = hphy_inst_PHYDDIODQOE_bus[25];
assign \phy_ddio_dqoe[26]  = hphy_inst_PHYDDIODQOE_bus[26];
assign \phy_ddio_dqoe[27]  = hphy_inst_PHYDDIODQOE_bus[27];
assign \phy_ddio_dqoe[28]  = hphy_inst_PHYDDIODQOE_bus[28];
assign \phy_ddio_dqoe[29]  = hphy_inst_PHYDDIODQOE_bus[29];
assign \phy_ddio_dqoe[30]  = hphy_inst_PHYDDIODQOE_bus[30];
assign \phy_ddio_dqoe[31]  = hphy_inst_PHYDDIODQOE_bus[31];
assign \phy_ddio_dqoe[32]  = hphy_inst_PHYDDIODQOE_bus[32];
assign \phy_ddio_dqoe[33]  = hphy_inst_PHYDDIODQOE_bus[33];
assign \phy_ddio_dqoe[36]  = hphy_inst_PHYDDIODQOE_bus[36];
assign \phy_ddio_dqoe[37]  = hphy_inst_PHYDDIODQOE_bus[37];
assign \phy_ddio_dqoe[38]  = hphy_inst_PHYDDIODQOE_bus[38];
assign \phy_ddio_dqoe[39]  = hphy_inst_PHYDDIODQOE_bus[39];
assign \phy_ddio_dqoe[40]  = hphy_inst_PHYDDIODQOE_bus[40];
assign \phy_ddio_dqoe[41]  = hphy_inst_PHYDDIODQOE_bus[41];
assign \phy_ddio_dqoe[42]  = hphy_inst_PHYDDIODQOE_bus[42];
assign \phy_ddio_dqoe[43]  = hphy_inst_PHYDDIODQOE_bus[43];
assign \phy_ddio_dqoe[44]  = hphy_inst_PHYDDIODQOE_bus[44];
assign \phy_ddio_dqoe[45]  = hphy_inst_PHYDDIODQOE_bus[45];
assign \phy_ddio_dqoe[46]  = hphy_inst_PHYDDIODQOE_bus[46];
assign \phy_ddio_dqoe[47]  = hphy_inst_PHYDDIODQOE_bus[47];
assign \phy_ddio_dqoe[48]  = hphy_inst_PHYDDIODQOE_bus[48];
assign \phy_ddio_dqoe[49]  = hphy_inst_PHYDDIODQOE_bus[49];
assign \phy_ddio_dqoe[50]  = hphy_inst_PHYDDIODQOE_bus[50];
assign \phy_ddio_dqoe[51]  = hphy_inst_PHYDDIODQOE_bus[51];
assign \phy_ddio_dqoe[54]  = hphy_inst_PHYDDIODQOE_bus[54];
assign \phy_ddio_dqoe[55]  = hphy_inst_PHYDDIODQOE_bus[55];
assign \phy_ddio_dqoe[56]  = hphy_inst_PHYDDIODQOE_bus[56];
assign \phy_ddio_dqoe[57]  = hphy_inst_PHYDDIODQOE_bus[57];
assign \phy_ddio_dqoe[58]  = hphy_inst_PHYDDIODQOE_bus[58];
assign \phy_ddio_dqoe[59]  = hphy_inst_PHYDDIODQOE_bus[59];
assign \phy_ddio_dqoe[60]  = hphy_inst_PHYDDIODQOE_bus[60];
assign \phy_ddio_dqoe[61]  = hphy_inst_PHYDDIODQOE_bus[61];
assign \phy_ddio_dqoe[62]  = hphy_inst_PHYDDIODQOE_bus[62];
assign \phy_ddio_dqoe[63]  = hphy_inst_PHYDDIODQOE_bus[63];
assign \phy_ddio_dqoe[64]  = hphy_inst_PHYDDIODQOE_bus[64];
assign \phy_ddio_dqoe[65]  = hphy_inst_PHYDDIODQOE_bus[65];
assign \phy_ddio_dqoe[66]  = hphy_inst_PHYDDIODQOE_bus[66];
assign \phy_ddio_dqoe[67]  = hphy_inst_PHYDDIODQOE_bus[67];
assign \phy_ddio_dqoe[68]  = hphy_inst_PHYDDIODQOE_bus[68];
assign \phy_ddio_dqoe[69]  = hphy_inst_PHYDDIODQOE_bus[69];

assign \phy_ddio_dqs_dout[0]  = hphy_inst_PHYDDIODQSDOUT_bus[0];
assign \phy_ddio_dqs_dout[1]  = hphy_inst_PHYDDIODQSDOUT_bus[1];
assign \phy_ddio_dqs_dout[2]  = hphy_inst_PHYDDIODQSDOUT_bus[2];
assign \phy_ddio_dqs_dout[3]  = hphy_inst_PHYDDIODQSDOUT_bus[3];
assign \phy_ddio_dqs_dout[4]  = hphy_inst_PHYDDIODQSDOUT_bus[4];
assign \phy_ddio_dqs_dout[5]  = hphy_inst_PHYDDIODQSDOUT_bus[5];
assign \phy_ddio_dqs_dout[6]  = hphy_inst_PHYDDIODQSDOUT_bus[6];
assign \phy_ddio_dqs_dout[7]  = hphy_inst_PHYDDIODQSDOUT_bus[7];
assign \phy_ddio_dqs_dout[8]  = hphy_inst_PHYDDIODQSDOUT_bus[8];
assign \phy_ddio_dqs_dout[9]  = hphy_inst_PHYDDIODQSDOUT_bus[9];
assign \phy_ddio_dqs_dout[10]  = hphy_inst_PHYDDIODQSDOUT_bus[10];
assign \phy_ddio_dqs_dout[11]  = hphy_inst_PHYDDIODQSDOUT_bus[11];
assign \phy_ddio_dqs_dout[12]  = hphy_inst_PHYDDIODQSDOUT_bus[12];
assign \phy_ddio_dqs_dout[13]  = hphy_inst_PHYDDIODQSDOUT_bus[13];
assign \phy_ddio_dqs_dout[14]  = hphy_inst_PHYDDIODQSDOUT_bus[14];
assign \phy_ddio_dqs_dout[15]  = hphy_inst_PHYDDIODQSDOUT_bus[15];

assign \phy_ddio_dqslogic_aclr_fifoctrl[0]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[0];
assign \phy_ddio_dqslogic_aclr_fifoctrl[1]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[1];
assign \phy_ddio_dqslogic_aclr_fifoctrl[2]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[2];
assign \phy_ddio_dqslogic_aclr_fifoctrl[3]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[3];

assign \phy_ddio_dqslogic_aclr_pstamble[0]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[0];
assign \phy_ddio_dqslogic_aclr_pstamble[1]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[1];
assign \phy_ddio_dqslogic_aclr_pstamble[2]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[2];
assign \phy_ddio_dqslogic_aclr_pstamble[3]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[3];

assign \phy_ddio_dqslogic_dqsena[0]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[0];
assign \phy_ddio_dqslogic_dqsena[1]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[1];
assign \phy_ddio_dqslogic_dqsena[2]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[2];
assign \phy_ddio_dqslogic_dqsena[3]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[3];
assign \phy_ddio_dqslogic_dqsena[4]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[4];
assign \phy_ddio_dqslogic_dqsena[5]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[5];
assign \phy_ddio_dqslogic_dqsena[6]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[6];
assign \phy_ddio_dqslogic_dqsena[7]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[7];

assign \phy_ddio_dqslogic_fiforeset[0]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[0];
assign \phy_ddio_dqslogic_fiforeset[1]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[1];
assign \phy_ddio_dqslogic_fiforeset[2]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[2];
assign \phy_ddio_dqslogic_fiforeset[3]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[3];

assign \phy_ddio_dqslogic_incrdataen[0]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[0];
assign \phy_ddio_dqslogic_incrdataen[1]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[1];
assign \phy_ddio_dqslogic_incrdataen[2]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[2];
assign \phy_ddio_dqslogic_incrdataen[3]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[3];
assign \phy_ddio_dqslogic_incrdataen[4]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[4];
assign \phy_ddio_dqslogic_incrdataen[5]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[5];
assign \phy_ddio_dqslogic_incrdataen[6]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[6];
assign \phy_ddio_dqslogic_incrdataen[7]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[7];

assign \phy_ddio_dqslogic_incwrptr[0]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[0];
assign \phy_ddio_dqslogic_incwrptr[1]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[1];
assign \phy_ddio_dqslogic_incwrptr[2]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[2];
assign \phy_ddio_dqslogic_incwrptr[3]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[3];
assign \phy_ddio_dqslogic_incwrptr[4]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[4];
assign \phy_ddio_dqslogic_incwrptr[5]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[5];
assign \phy_ddio_dqslogic_incwrptr[6]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[6];
assign \phy_ddio_dqslogic_incwrptr[7]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[7];

assign \phy_ddio_dqslogic_oct[0]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[0];
assign \phy_ddio_dqslogic_oct[1]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[1];
assign \phy_ddio_dqslogic_oct[2]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[2];
assign \phy_ddio_dqslogic_oct[3]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[3];
assign \phy_ddio_dqslogic_oct[4]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[4];
assign \phy_ddio_dqslogic_oct[5]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[5];
assign \phy_ddio_dqslogic_oct[6]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[6];
assign \phy_ddio_dqslogic_oct[7]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[7];

assign \phy_ddio_dqslogic_readlatency[0]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[0];
assign \phy_ddio_dqslogic_readlatency[1]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[1];
assign \phy_ddio_dqslogic_readlatency[2]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[2];
assign \phy_ddio_dqslogic_readlatency[3]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[3];
assign \phy_ddio_dqslogic_readlatency[4]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[4];
assign \phy_ddio_dqslogic_readlatency[5]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[5];
assign \phy_ddio_dqslogic_readlatency[6]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[6];
assign \phy_ddio_dqslogic_readlatency[7]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[7];
assign \phy_ddio_dqslogic_readlatency[8]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[8];
assign \phy_ddio_dqslogic_readlatency[9]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[9];
assign \phy_ddio_dqslogic_readlatency[10]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[10];
assign \phy_ddio_dqslogic_readlatency[11]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[11];
assign \phy_ddio_dqslogic_readlatency[12]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[12];
assign \phy_ddio_dqslogic_readlatency[13]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[13];
assign \phy_ddio_dqslogic_readlatency[14]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[14];
assign \phy_ddio_dqslogic_readlatency[15]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[15];
assign \phy_ddio_dqslogic_readlatency[16]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[16];
assign \phy_ddio_dqslogic_readlatency[17]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[17];
assign \phy_ddio_dqslogic_readlatency[18]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[18];
assign \phy_ddio_dqslogic_readlatency[19]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[19];

assign \phy_ddio_dqs_oe[0]  = hphy_inst_PHYDDIODQSOE_bus[0];
assign \phy_ddio_dqs_oe[1]  = hphy_inst_PHYDDIODQSOE_bus[1];
assign \phy_ddio_dqs_oe[2]  = hphy_inst_PHYDDIODQSOE_bus[2];
assign \phy_ddio_dqs_oe[3]  = hphy_inst_PHYDDIODQSOE_bus[3];
assign \phy_ddio_dqs_oe[4]  = hphy_inst_PHYDDIODQSOE_bus[4];
assign \phy_ddio_dqs_oe[5]  = hphy_inst_PHYDDIODQSOE_bus[5];
assign \phy_ddio_dqs_oe[6]  = hphy_inst_PHYDDIODQSOE_bus[6];
assign \phy_ddio_dqs_oe[7]  = hphy_inst_PHYDDIODQSOE_bus[7];

assign \phy_ddio_odt[0]  = hphy_inst_PHYDDIOODTDOUT_bus[0];
assign \phy_ddio_odt[1]  = hphy_inst_PHYDDIOODTDOUT_bus[1];
assign \phy_ddio_odt[2]  = hphy_inst_PHYDDIOODTDOUT_bus[2];
assign \phy_ddio_odt[3]  = hphy_inst_PHYDDIOODTDOUT_bus[3];

assign \phy_ddio_ras_n[0]  = hphy_inst_PHYDDIORASNDOUT_bus[0];
assign \phy_ddio_ras_n[1]  = hphy_inst_PHYDDIORASNDOUT_bus[1];
assign \phy_ddio_ras_n[2]  = hphy_inst_PHYDDIORASNDOUT_bus[2];
assign \phy_ddio_ras_n[3]  = hphy_inst_PHYDDIORASNDOUT_bus[3];

assign \phy_ddio_reset_n[0]  = hphy_inst_PHYDDIORESETNDOUT_bus[0];
assign \phy_ddio_reset_n[1]  = hphy_inst_PHYDDIORESETNDOUT_bus[1];
assign \phy_ddio_reset_n[2]  = hphy_inst_PHYDDIORESETNDOUT_bus[2];
assign \phy_ddio_reset_n[3]  = hphy_inst_PHYDDIORESETNDOUT_bus[3];

assign \phy_ddio_we_n[0]  = hphy_inst_PHYDDIOWENDOUT_bus[0];
assign \phy_ddio_we_n[1]  = hphy_inst_PHYDDIOWENDOUT_bus[1];
assign \phy_ddio_we_n[2]  = hphy_inst_PHYDDIOWENDOUT_bus[2];
assign \phy_ddio_we_n[3]  = hphy_inst_PHYDDIOWENDOUT_bus[3];

Computer_System_hps_sdram_p0_acv_hard_io_pads uio_pads(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(\phy_ddio_address[0] ),
	.phy_ddio_address_1(\phy_ddio_address[1] ),
	.phy_ddio_address_2(\phy_ddio_address[2] ),
	.phy_ddio_address_3(\phy_ddio_address[3] ),
	.phy_ddio_address_4(\phy_ddio_address[4] ),
	.phy_ddio_address_5(\phy_ddio_address[5] ),
	.phy_ddio_address_6(\phy_ddio_address[6] ),
	.phy_ddio_address_7(\phy_ddio_address[7] ),
	.phy_ddio_address_8(\phy_ddio_address[8] ),
	.phy_ddio_address_9(\phy_ddio_address[9] ),
	.phy_ddio_address_10(\phy_ddio_address[10] ),
	.phy_ddio_address_11(\phy_ddio_address[11] ),
	.phy_ddio_address_12(\phy_ddio_address[12] ),
	.phy_ddio_address_13(\phy_ddio_address[13] ),
	.phy_ddio_address_14(\phy_ddio_address[14] ),
	.phy_ddio_address_15(\phy_ddio_address[15] ),
	.phy_ddio_address_16(\phy_ddio_address[16] ),
	.phy_ddio_address_17(\phy_ddio_address[17] ),
	.phy_ddio_address_18(\phy_ddio_address[18] ),
	.phy_ddio_address_19(\phy_ddio_address[19] ),
	.phy_ddio_address_20(\phy_ddio_address[20] ),
	.phy_ddio_address_21(\phy_ddio_address[21] ),
	.phy_ddio_address_22(\phy_ddio_address[22] ),
	.phy_ddio_address_23(\phy_ddio_address[23] ),
	.phy_ddio_address_24(\phy_ddio_address[24] ),
	.phy_ddio_address_25(\phy_ddio_address[25] ),
	.phy_ddio_address_26(\phy_ddio_address[26] ),
	.phy_ddio_address_27(\phy_ddio_address[27] ),
	.phy_ddio_address_28(\phy_ddio_address[28] ),
	.phy_ddio_address_29(\phy_ddio_address[29] ),
	.phy_ddio_address_30(\phy_ddio_address[30] ),
	.phy_ddio_address_31(\phy_ddio_address[31] ),
	.phy_ddio_address_32(\phy_ddio_address[32] ),
	.phy_ddio_address_33(\phy_ddio_address[33] ),
	.phy_ddio_address_34(\phy_ddio_address[34] ),
	.phy_ddio_address_35(\phy_ddio_address[35] ),
	.phy_ddio_address_36(\phy_ddio_address[36] ),
	.phy_ddio_address_37(\phy_ddio_address[37] ),
	.phy_ddio_address_38(\phy_ddio_address[38] ),
	.phy_ddio_address_39(\phy_ddio_address[39] ),
	.phy_ddio_address_40(\phy_ddio_address[40] ),
	.phy_ddio_address_41(\phy_ddio_address[41] ),
	.phy_ddio_address_42(\phy_ddio_address[42] ),
	.phy_ddio_address_43(\phy_ddio_address[43] ),
	.phy_ddio_address_44(\phy_ddio_address[44] ),
	.phy_ddio_address_45(\phy_ddio_address[45] ),
	.phy_ddio_address_46(\phy_ddio_address[46] ),
	.phy_ddio_address_47(\phy_ddio_address[47] ),
	.phy_ddio_address_48(\phy_ddio_address[48] ),
	.phy_ddio_address_49(\phy_ddio_address[49] ),
	.phy_ddio_address_50(\phy_ddio_address[50] ),
	.phy_ddio_address_51(\phy_ddio_address[51] ),
	.phy_ddio_address_52(\phy_ddio_address[52] ),
	.phy_ddio_address_53(\phy_ddio_address[53] ),
	.phy_ddio_address_54(\phy_ddio_address[54] ),
	.phy_ddio_address_55(\phy_ddio_address[55] ),
	.phy_ddio_address_56(\phy_ddio_address[56] ),
	.phy_ddio_address_57(\phy_ddio_address[57] ),
	.phy_ddio_address_58(\phy_ddio_address[58] ),
	.phy_ddio_address_59(\phy_ddio_address[59] ),
	.phy_ddio_bank_0(\phy_ddio_bank[0] ),
	.phy_ddio_bank_1(\phy_ddio_bank[1] ),
	.phy_ddio_bank_2(\phy_ddio_bank[2] ),
	.phy_ddio_bank_3(\phy_ddio_bank[3] ),
	.phy_ddio_bank_4(\phy_ddio_bank[4] ),
	.phy_ddio_bank_5(\phy_ddio_bank[5] ),
	.phy_ddio_bank_6(\phy_ddio_bank[6] ),
	.phy_ddio_bank_7(\phy_ddio_bank[7] ),
	.phy_ddio_bank_8(\phy_ddio_bank[8] ),
	.phy_ddio_bank_9(\phy_ddio_bank[9] ),
	.phy_ddio_bank_10(\phy_ddio_bank[10] ),
	.phy_ddio_bank_11(\phy_ddio_bank[11] ),
	.phy_ddio_cas_n_0(\phy_ddio_cas_n[0] ),
	.phy_ddio_cas_n_1(\phy_ddio_cas_n[1] ),
	.phy_ddio_cas_n_2(\phy_ddio_cas_n[2] ),
	.phy_ddio_cas_n_3(\phy_ddio_cas_n[3] ),
	.phy_ddio_ck_0(\phy_ddio_ck[0] ),
	.phy_ddio_ck_1(\phy_ddio_ck[1] ),
	.phy_ddio_cke_0(\phy_ddio_cke[0] ),
	.phy_ddio_cke_1(\phy_ddio_cke[1] ),
	.phy_ddio_cke_2(\phy_ddio_cke[2] ),
	.phy_ddio_cke_3(\phy_ddio_cke[3] ),
	.phy_ddio_cs_n_0(\phy_ddio_cs_n[0] ),
	.phy_ddio_cs_n_1(\phy_ddio_cs_n[1] ),
	.phy_ddio_cs_n_2(\phy_ddio_cs_n[2] ),
	.phy_ddio_cs_n_3(\phy_ddio_cs_n[3] ),
	.phy_ddio_dmdout_0(\phy_ddio_dmdout[0] ),
	.phy_ddio_dmdout_1(\phy_ddio_dmdout[1] ),
	.phy_ddio_dmdout_2(\phy_ddio_dmdout[2] ),
	.phy_ddio_dmdout_3(\phy_ddio_dmdout[3] ),
	.phy_ddio_dmdout_4(\phy_ddio_dmdout[4] ),
	.phy_ddio_dmdout_5(\phy_ddio_dmdout[5] ),
	.phy_ddio_dmdout_6(\phy_ddio_dmdout[6] ),
	.phy_ddio_dmdout_7(\phy_ddio_dmdout[7] ),
	.phy_ddio_dmdout_8(\phy_ddio_dmdout[8] ),
	.phy_ddio_dmdout_9(\phy_ddio_dmdout[9] ),
	.phy_ddio_dmdout_10(\phy_ddio_dmdout[10] ),
	.phy_ddio_dmdout_11(\phy_ddio_dmdout[11] ),
	.phy_ddio_dmdout_12(\phy_ddio_dmdout[12] ),
	.phy_ddio_dmdout_13(\phy_ddio_dmdout[13] ),
	.phy_ddio_dmdout_14(\phy_ddio_dmdout[14] ),
	.phy_ddio_dmdout_15(\phy_ddio_dmdout[15] ),
	.phy_ddio_dqdout_0(\phy_ddio_dqdout[0] ),
	.phy_ddio_dqdout_1(\phy_ddio_dqdout[1] ),
	.phy_ddio_dqdout_2(\phy_ddio_dqdout[2] ),
	.phy_ddio_dqdout_3(\phy_ddio_dqdout[3] ),
	.phy_ddio_dqdout_4(\phy_ddio_dqdout[4] ),
	.phy_ddio_dqdout_5(\phy_ddio_dqdout[5] ),
	.phy_ddio_dqdout_6(\phy_ddio_dqdout[6] ),
	.phy_ddio_dqdout_7(\phy_ddio_dqdout[7] ),
	.phy_ddio_dqdout_8(\phy_ddio_dqdout[8] ),
	.phy_ddio_dqdout_9(\phy_ddio_dqdout[9] ),
	.phy_ddio_dqdout_10(\phy_ddio_dqdout[10] ),
	.phy_ddio_dqdout_11(\phy_ddio_dqdout[11] ),
	.phy_ddio_dqdout_12(\phy_ddio_dqdout[12] ),
	.phy_ddio_dqdout_13(\phy_ddio_dqdout[13] ),
	.phy_ddio_dqdout_14(\phy_ddio_dqdout[14] ),
	.phy_ddio_dqdout_15(\phy_ddio_dqdout[15] ),
	.phy_ddio_dqdout_16(\phy_ddio_dqdout[16] ),
	.phy_ddio_dqdout_17(\phy_ddio_dqdout[17] ),
	.phy_ddio_dqdout_18(\phy_ddio_dqdout[18] ),
	.phy_ddio_dqdout_19(\phy_ddio_dqdout[19] ),
	.phy_ddio_dqdout_20(\phy_ddio_dqdout[20] ),
	.phy_ddio_dqdout_21(\phy_ddio_dqdout[21] ),
	.phy_ddio_dqdout_22(\phy_ddio_dqdout[22] ),
	.phy_ddio_dqdout_23(\phy_ddio_dqdout[23] ),
	.phy_ddio_dqdout_24(\phy_ddio_dqdout[24] ),
	.phy_ddio_dqdout_25(\phy_ddio_dqdout[25] ),
	.phy_ddio_dqdout_26(\phy_ddio_dqdout[26] ),
	.phy_ddio_dqdout_27(\phy_ddio_dqdout[27] ),
	.phy_ddio_dqdout_28(\phy_ddio_dqdout[28] ),
	.phy_ddio_dqdout_29(\phy_ddio_dqdout[29] ),
	.phy_ddio_dqdout_30(\phy_ddio_dqdout[30] ),
	.phy_ddio_dqdout_31(\phy_ddio_dqdout[31] ),
	.phy_ddio_dqdout_36(\phy_ddio_dqdout[36] ),
	.phy_ddio_dqdout_37(\phy_ddio_dqdout[37] ),
	.phy_ddio_dqdout_38(\phy_ddio_dqdout[38] ),
	.phy_ddio_dqdout_39(\phy_ddio_dqdout[39] ),
	.phy_ddio_dqdout_40(\phy_ddio_dqdout[40] ),
	.phy_ddio_dqdout_41(\phy_ddio_dqdout[41] ),
	.phy_ddio_dqdout_42(\phy_ddio_dqdout[42] ),
	.phy_ddio_dqdout_43(\phy_ddio_dqdout[43] ),
	.phy_ddio_dqdout_44(\phy_ddio_dqdout[44] ),
	.phy_ddio_dqdout_45(\phy_ddio_dqdout[45] ),
	.phy_ddio_dqdout_46(\phy_ddio_dqdout[46] ),
	.phy_ddio_dqdout_47(\phy_ddio_dqdout[47] ),
	.phy_ddio_dqdout_48(\phy_ddio_dqdout[48] ),
	.phy_ddio_dqdout_49(\phy_ddio_dqdout[49] ),
	.phy_ddio_dqdout_50(\phy_ddio_dqdout[50] ),
	.phy_ddio_dqdout_51(\phy_ddio_dqdout[51] ),
	.phy_ddio_dqdout_52(\phy_ddio_dqdout[52] ),
	.phy_ddio_dqdout_53(\phy_ddio_dqdout[53] ),
	.phy_ddio_dqdout_54(\phy_ddio_dqdout[54] ),
	.phy_ddio_dqdout_55(\phy_ddio_dqdout[55] ),
	.phy_ddio_dqdout_56(\phy_ddio_dqdout[56] ),
	.phy_ddio_dqdout_57(\phy_ddio_dqdout[57] ),
	.phy_ddio_dqdout_58(\phy_ddio_dqdout[58] ),
	.phy_ddio_dqdout_59(\phy_ddio_dqdout[59] ),
	.phy_ddio_dqdout_60(\phy_ddio_dqdout[60] ),
	.phy_ddio_dqdout_61(\phy_ddio_dqdout[61] ),
	.phy_ddio_dqdout_62(\phy_ddio_dqdout[62] ),
	.phy_ddio_dqdout_63(\phy_ddio_dqdout[63] ),
	.phy_ddio_dqdout_64(\phy_ddio_dqdout[64] ),
	.phy_ddio_dqdout_65(\phy_ddio_dqdout[65] ),
	.phy_ddio_dqdout_66(\phy_ddio_dqdout[66] ),
	.phy_ddio_dqdout_67(\phy_ddio_dqdout[67] ),
	.phy_ddio_dqdout_72(\phy_ddio_dqdout[72] ),
	.phy_ddio_dqdout_73(\phy_ddio_dqdout[73] ),
	.phy_ddio_dqdout_74(\phy_ddio_dqdout[74] ),
	.phy_ddio_dqdout_75(\phy_ddio_dqdout[75] ),
	.phy_ddio_dqdout_76(\phy_ddio_dqdout[76] ),
	.phy_ddio_dqdout_77(\phy_ddio_dqdout[77] ),
	.phy_ddio_dqdout_78(\phy_ddio_dqdout[78] ),
	.phy_ddio_dqdout_79(\phy_ddio_dqdout[79] ),
	.phy_ddio_dqdout_80(\phy_ddio_dqdout[80] ),
	.phy_ddio_dqdout_81(\phy_ddio_dqdout[81] ),
	.phy_ddio_dqdout_82(\phy_ddio_dqdout[82] ),
	.phy_ddio_dqdout_83(\phy_ddio_dqdout[83] ),
	.phy_ddio_dqdout_84(\phy_ddio_dqdout[84] ),
	.phy_ddio_dqdout_85(\phy_ddio_dqdout[85] ),
	.phy_ddio_dqdout_86(\phy_ddio_dqdout[86] ),
	.phy_ddio_dqdout_87(\phy_ddio_dqdout[87] ),
	.phy_ddio_dqdout_88(\phy_ddio_dqdout[88] ),
	.phy_ddio_dqdout_89(\phy_ddio_dqdout[89] ),
	.phy_ddio_dqdout_90(\phy_ddio_dqdout[90] ),
	.phy_ddio_dqdout_91(\phy_ddio_dqdout[91] ),
	.phy_ddio_dqdout_92(\phy_ddio_dqdout[92] ),
	.phy_ddio_dqdout_93(\phy_ddio_dqdout[93] ),
	.phy_ddio_dqdout_94(\phy_ddio_dqdout[94] ),
	.phy_ddio_dqdout_95(\phy_ddio_dqdout[95] ),
	.phy_ddio_dqdout_96(\phy_ddio_dqdout[96] ),
	.phy_ddio_dqdout_97(\phy_ddio_dqdout[97] ),
	.phy_ddio_dqdout_98(\phy_ddio_dqdout[98] ),
	.phy_ddio_dqdout_99(\phy_ddio_dqdout[99] ),
	.phy_ddio_dqdout_100(\phy_ddio_dqdout[100] ),
	.phy_ddio_dqdout_101(\phy_ddio_dqdout[101] ),
	.phy_ddio_dqdout_102(\phy_ddio_dqdout[102] ),
	.phy_ddio_dqdout_103(\phy_ddio_dqdout[103] ),
	.phy_ddio_dqdout_108(\phy_ddio_dqdout[108] ),
	.phy_ddio_dqdout_109(\phy_ddio_dqdout[109] ),
	.phy_ddio_dqdout_110(\phy_ddio_dqdout[110] ),
	.phy_ddio_dqdout_111(\phy_ddio_dqdout[111] ),
	.phy_ddio_dqdout_112(\phy_ddio_dqdout[112] ),
	.phy_ddio_dqdout_113(\phy_ddio_dqdout[113] ),
	.phy_ddio_dqdout_114(\phy_ddio_dqdout[114] ),
	.phy_ddio_dqdout_115(\phy_ddio_dqdout[115] ),
	.phy_ddio_dqdout_116(\phy_ddio_dqdout[116] ),
	.phy_ddio_dqdout_117(\phy_ddio_dqdout[117] ),
	.phy_ddio_dqdout_118(\phy_ddio_dqdout[118] ),
	.phy_ddio_dqdout_119(\phy_ddio_dqdout[119] ),
	.phy_ddio_dqdout_120(\phy_ddio_dqdout[120] ),
	.phy_ddio_dqdout_121(\phy_ddio_dqdout[121] ),
	.phy_ddio_dqdout_122(\phy_ddio_dqdout[122] ),
	.phy_ddio_dqdout_123(\phy_ddio_dqdout[123] ),
	.phy_ddio_dqdout_124(\phy_ddio_dqdout[124] ),
	.phy_ddio_dqdout_125(\phy_ddio_dqdout[125] ),
	.phy_ddio_dqdout_126(\phy_ddio_dqdout[126] ),
	.phy_ddio_dqdout_127(\phy_ddio_dqdout[127] ),
	.phy_ddio_dqdout_128(\phy_ddio_dqdout[128] ),
	.phy_ddio_dqdout_129(\phy_ddio_dqdout[129] ),
	.phy_ddio_dqdout_130(\phy_ddio_dqdout[130] ),
	.phy_ddio_dqdout_131(\phy_ddio_dqdout[131] ),
	.phy_ddio_dqdout_132(\phy_ddio_dqdout[132] ),
	.phy_ddio_dqdout_133(\phy_ddio_dqdout[133] ),
	.phy_ddio_dqdout_134(\phy_ddio_dqdout[134] ),
	.phy_ddio_dqdout_135(\phy_ddio_dqdout[135] ),
	.phy_ddio_dqdout_136(\phy_ddio_dqdout[136] ),
	.phy_ddio_dqdout_137(\phy_ddio_dqdout[137] ),
	.phy_ddio_dqdout_138(\phy_ddio_dqdout[138] ),
	.phy_ddio_dqdout_139(\phy_ddio_dqdout[139] ),
	.phy_ddio_dqoe_0(\phy_ddio_dqoe[0] ),
	.phy_ddio_dqoe_1(\phy_ddio_dqoe[1] ),
	.phy_ddio_dqoe_2(\phy_ddio_dqoe[2] ),
	.phy_ddio_dqoe_3(\phy_ddio_dqoe[3] ),
	.phy_ddio_dqoe_4(\phy_ddio_dqoe[4] ),
	.phy_ddio_dqoe_5(\phy_ddio_dqoe[5] ),
	.phy_ddio_dqoe_6(\phy_ddio_dqoe[6] ),
	.phy_ddio_dqoe_7(\phy_ddio_dqoe[7] ),
	.phy_ddio_dqoe_8(\phy_ddio_dqoe[8] ),
	.phy_ddio_dqoe_9(\phy_ddio_dqoe[9] ),
	.phy_ddio_dqoe_10(\phy_ddio_dqoe[10] ),
	.phy_ddio_dqoe_11(\phy_ddio_dqoe[11] ),
	.phy_ddio_dqoe_12(\phy_ddio_dqoe[12] ),
	.phy_ddio_dqoe_13(\phy_ddio_dqoe[13] ),
	.phy_ddio_dqoe_14(\phy_ddio_dqoe[14] ),
	.phy_ddio_dqoe_15(\phy_ddio_dqoe[15] ),
	.phy_ddio_dqoe_18(\phy_ddio_dqoe[18] ),
	.phy_ddio_dqoe_19(\phy_ddio_dqoe[19] ),
	.phy_ddio_dqoe_20(\phy_ddio_dqoe[20] ),
	.phy_ddio_dqoe_21(\phy_ddio_dqoe[21] ),
	.phy_ddio_dqoe_22(\phy_ddio_dqoe[22] ),
	.phy_ddio_dqoe_23(\phy_ddio_dqoe[23] ),
	.phy_ddio_dqoe_24(\phy_ddio_dqoe[24] ),
	.phy_ddio_dqoe_25(\phy_ddio_dqoe[25] ),
	.phy_ddio_dqoe_26(\phy_ddio_dqoe[26] ),
	.phy_ddio_dqoe_27(\phy_ddio_dqoe[27] ),
	.phy_ddio_dqoe_28(\phy_ddio_dqoe[28] ),
	.phy_ddio_dqoe_29(\phy_ddio_dqoe[29] ),
	.phy_ddio_dqoe_30(\phy_ddio_dqoe[30] ),
	.phy_ddio_dqoe_31(\phy_ddio_dqoe[31] ),
	.phy_ddio_dqoe_32(\phy_ddio_dqoe[32] ),
	.phy_ddio_dqoe_33(\phy_ddio_dqoe[33] ),
	.phy_ddio_dqoe_36(\phy_ddio_dqoe[36] ),
	.phy_ddio_dqoe_37(\phy_ddio_dqoe[37] ),
	.phy_ddio_dqoe_38(\phy_ddio_dqoe[38] ),
	.phy_ddio_dqoe_39(\phy_ddio_dqoe[39] ),
	.phy_ddio_dqoe_40(\phy_ddio_dqoe[40] ),
	.phy_ddio_dqoe_41(\phy_ddio_dqoe[41] ),
	.phy_ddio_dqoe_42(\phy_ddio_dqoe[42] ),
	.phy_ddio_dqoe_43(\phy_ddio_dqoe[43] ),
	.phy_ddio_dqoe_44(\phy_ddio_dqoe[44] ),
	.phy_ddio_dqoe_45(\phy_ddio_dqoe[45] ),
	.phy_ddio_dqoe_46(\phy_ddio_dqoe[46] ),
	.phy_ddio_dqoe_47(\phy_ddio_dqoe[47] ),
	.phy_ddio_dqoe_48(\phy_ddio_dqoe[48] ),
	.phy_ddio_dqoe_49(\phy_ddio_dqoe[49] ),
	.phy_ddio_dqoe_50(\phy_ddio_dqoe[50] ),
	.phy_ddio_dqoe_51(\phy_ddio_dqoe[51] ),
	.phy_ddio_dqoe_54(\phy_ddio_dqoe[54] ),
	.phy_ddio_dqoe_55(\phy_ddio_dqoe[55] ),
	.phy_ddio_dqoe_56(\phy_ddio_dqoe[56] ),
	.phy_ddio_dqoe_57(\phy_ddio_dqoe[57] ),
	.phy_ddio_dqoe_58(\phy_ddio_dqoe[58] ),
	.phy_ddio_dqoe_59(\phy_ddio_dqoe[59] ),
	.phy_ddio_dqoe_60(\phy_ddio_dqoe[60] ),
	.phy_ddio_dqoe_61(\phy_ddio_dqoe[61] ),
	.phy_ddio_dqoe_62(\phy_ddio_dqoe[62] ),
	.phy_ddio_dqoe_63(\phy_ddio_dqoe[63] ),
	.phy_ddio_dqoe_64(\phy_ddio_dqoe[64] ),
	.phy_ddio_dqoe_65(\phy_ddio_dqoe[65] ),
	.phy_ddio_dqoe_66(\phy_ddio_dqoe[66] ),
	.phy_ddio_dqoe_67(\phy_ddio_dqoe[67] ),
	.phy_ddio_dqoe_68(\phy_ddio_dqoe[68] ),
	.phy_ddio_dqoe_69(\phy_ddio_dqoe[69] ),
	.phy_ddio_dqs_dout_0(\phy_ddio_dqs_dout[0] ),
	.phy_ddio_dqs_dout_1(\phy_ddio_dqs_dout[1] ),
	.phy_ddio_dqs_dout_2(\phy_ddio_dqs_dout[2] ),
	.phy_ddio_dqs_dout_3(\phy_ddio_dqs_dout[3] ),
	.phy_ddio_dqs_dout_4(\phy_ddio_dqs_dout[4] ),
	.phy_ddio_dqs_dout_5(\phy_ddio_dqs_dout[5] ),
	.phy_ddio_dqs_dout_6(\phy_ddio_dqs_dout[6] ),
	.phy_ddio_dqs_dout_7(\phy_ddio_dqs_dout[7] ),
	.phy_ddio_dqs_dout_8(\phy_ddio_dqs_dout[8] ),
	.phy_ddio_dqs_dout_9(\phy_ddio_dqs_dout[9] ),
	.phy_ddio_dqs_dout_10(\phy_ddio_dqs_dout[10] ),
	.phy_ddio_dqs_dout_11(\phy_ddio_dqs_dout[11] ),
	.phy_ddio_dqs_dout_12(\phy_ddio_dqs_dout[12] ),
	.phy_ddio_dqs_dout_13(\phy_ddio_dqs_dout[13] ),
	.phy_ddio_dqs_dout_14(\phy_ddio_dqs_dout[14] ),
	.phy_ddio_dqs_dout_15(\phy_ddio_dqs_dout[15] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(\phy_ddio_dqslogic_aclr_fifoctrl[0] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(\phy_ddio_dqslogic_aclr_fifoctrl[1] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(\phy_ddio_dqslogic_aclr_fifoctrl[2] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(\phy_ddio_dqslogic_aclr_fifoctrl[3] ),
	.phy_ddio_dqslogic_aclr_pstamble_0(\phy_ddio_dqslogic_aclr_pstamble[0] ),
	.phy_ddio_dqslogic_aclr_pstamble_1(\phy_ddio_dqslogic_aclr_pstamble[1] ),
	.phy_ddio_dqslogic_aclr_pstamble_2(\phy_ddio_dqslogic_aclr_pstamble[2] ),
	.phy_ddio_dqslogic_aclr_pstamble_3(\phy_ddio_dqslogic_aclr_pstamble[3] ),
	.phy_ddio_dqslogic_dqsena_0(\phy_ddio_dqslogic_dqsena[0] ),
	.phy_ddio_dqslogic_dqsena_1(\phy_ddio_dqslogic_dqsena[1] ),
	.phy_ddio_dqslogic_dqsena_2(\phy_ddio_dqslogic_dqsena[2] ),
	.phy_ddio_dqslogic_dqsena_3(\phy_ddio_dqslogic_dqsena[3] ),
	.phy_ddio_dqslogic_dqsena_4(\phy_ddio_dqslogic_dqsena[4] ),
	.phy_ddio_dqslogic_dqsena_5(\phy_ddio_dqslogic_dqsena[5] ),
	.phy_ddio_dqslogic_dqsena_6(\phy_ddio_dqslogic_dqsena[6] ),
	.phy_ddio_dqslogic_dqsena_7(\phy_ddio_dqslogic_dqsena[7] ),
	.phy_ddio_dqslogic_fiforeset_0(\phy_ddio_dqslogic_fiforeset[0] ),
	.phy_ddio_dqslogic_fiforeset_1(\phy_ddio_dqslogic_fiforeset[1] ),
	.phy_ddio_dqslogic_fiforeset_2(\phy_ddio_dqslogic_fiforeset[2] ),
	.phy_ddio_dqslogic_fiforeset_3(\phy_ddio_dqslogic_fiforeset[3] ),
	.phy_ddio_dqslogic_incrdataen_0(\phy_ddio_dqslogic_incrdataen[0] ),
	.phy_ddio_dqslogic_incrdataen_1(\phy_ddio_dqslogic_incrdataen[1] ),
	.phy_ddio_dqslogic_incrdataen_2(\phy_ddio_dqslogic_incrdataen[2] ),
	.phy_ddio_dqslogic_incrdataen_3(\phy_ddio_dqslogic_incrdataen[3] ),
	.phy_ddio_dqslogic_incrdataen_4(\phy_ddio_dqslogic_incrdataen[4] ),
	.phy_ddio_dqslogic_incrdataen_5(\phy_ddio_dqslogic_incrdataen[5] ),
	.phy_ddio_dqslogic_incrdataen_6(\phy_ddio_dqslogic_incrdataen[6] ),
	.phy_ddio_dqslogic_incrdataen_7(\phy_ddio_dqslogic_incrdataen[7] ),
	.phy_ddio_dqslogic_incwrptr_0(\phy_ddio_dqslogic_incwrptr[0] ),
	.phy_ddio_dqslogic_incwrptr_1(\phy_ddio_dqslogic_incwrptr[1] ),
	.phy_ddio_dqslogic_incwrptr_2(\phy_ddio_dqslogic_incwrptr[2] ),
	.phy_ddio_dqslogic_incwrptr_3(\phy_ddio_dqslogic_incwrptr[3] ),
	.phy_ddio_dqslogic_incwrptr_4(\phy_ddio_dqslogic_incwrptr[4] ),
	.phy_ddio_dqslogic_incwrptr_5(\phy_ddio_dqslogic_incwrptr[5] ),
	.phy_ddio_dqslogic_incwrptr_6(\phy_ddio_dqslogic_incwrptr[6] ),
	.phy_ddio_dqslogic_incwrptr_7(\phy_ddio_dqslogic_incwrptr[7] ),
	.phy_ddio_dqslogic_oct_0(\phy_ddio_dqslogic_oct[0] ),
	.phy_ddio_dqslogic_oct_1(\phy_ddio_dqslogic_oct[1] ),
	.phy_ddio_dqslogic_oct_2(\phy_ddio_dqslogic_oct[2] ),
	.phy_ddio_dqslogic_oct_3(\phy_ddio_dqslogic_oct[3] ),
	.phy_ddio_dqslogic_oct_4(\phy_ddio_dqslogic_oct[4] ),
	.phy_ddio_dqslogic_oct_5(\phy_ddio_dqslogic_oct[5] ),
	.phy_ddio_dqslogic_oct_6(\phy_ddio_dqslogic_oct[6] ),
	.phy_ddio_dqslogic_oct_7(\phy_ddio_dqslogic_oct[7] ),
	.phy_ddio_dqslogic_readlatency_0(\phy_ddio_dqslogic_readlatency[0] ),
	.phy_ddio_dqslogic_readlatency_1(\phy_ddio_dqslogic_readlatency[1] ),
	.phy_ddio_dqslogic_readlatency_2(\phy_ddio_dqslogic_readlatency[2] ),
	.phy_ddio_dqslogic_readlatency_3(\phy_ddio_dqslogic_readlatency[3] ),
	.phy_ddio_dqslogic_readlatency_4(\phy_ddio_dqslogic_readlatency[4] ),
	.phy_ddio_dqslogic_readlatency_5(\phy_ddio_dqslogic_readlatency[5] ),
	.phy_ddio_dqslogic_readlatency_6(\phy_ddio_dqslogic_readlatency[6] ),
	.phy_ddio_dqslogic_readlatency_7(\phy_ddio_dqslogic_readlatency[7] ),
	.phy_ddio_dqslogic_readlatency_8(\phy_ddio_dqslogic_readlatency[8] ),
	.phy_ddio_dqslogic_readlatency_9(\phy_ddio_dqslogic_readlatency[9] ),
	.phy_ddio_dqslogic_readlatency_10(\phy_ddio_dqslogic_readlatency[10] ),
	.phy_ddio_dqslogic_readlatency_11(\phy_ddio_dqslogic_readlatency[11] ),
	.phy_ddio_dqslogic_readlatency_12(\phy_ddio_dqslogic_readlatency[12] ),
	.phy_ddio_dqslogic_readlatency_13(\phy_ddio_dqslogic_readlatency[13] ),
	.phy_ddio_dqslogic_readlatency_14(\phy_ddio_dqslogic_readlatency[14] ),
	.phy_ddio_dqslogic_readlatency_15(\phy_ddio_dqslogic_readlatency[15] ),
	.phy_ddio_dqslogic_readlatency_16(\phy_ddio_dqslogic_readlatency[16] ),
	.phy_ddio_dqslogic_readlatency_17(\phy_ddio_dqslogic_readlatency[17] ),
	.phy_ddio_dqslogic_readlatency_18(\phy_ddio_dqslogic_readlatency[18] ),
	.phy_ddio_dqslogic_readlatency_19(\phy_ddio_dqslogic_readlatency[19] ),
	.phy_ddio_dqs_oe_0(\phy_ddio_dqs_oe[0] ),
	.phy_ddio_dqs_oe_1(\phy_ddio_dqs_oe[1] ),
	.phy_ddio_dqs_oe_2(\phy_ddio_dqs_oe[2] ),
	.phy_ddio_dqs_oe_3(\phy_ddio_dqs_oe[3] ),
	.phy_ddio_dqs_oe_4(\phy_ddio_dqs_oe[4] ),
	.phy_ddio_dqs_oe_5(\phy_ddio_dqs_oe[5] ),
	.phy_ddio_dqs_oe_6(\phy_ddio_dqs_oe[6] ),
	.phy_ddio_dqs_oe_7(\phy_ddio_dqs_oe[7] ),
	.phy_ddio_odt_0(\phy_ddio_odt[0] ),
	.phy_ddio_odt_1(\phy_ddio_odt[1] ),
	.phy_ddio_odt_2(\phy_ddio_odt[2] ),
	.phy_ddio_odt_3(\phy_ddio_odt[3] ),
	.phy_ddio_ras_n_0(\phy_ddio_ras_n[0] ),
	.phy_ddio_ras_n_1(\phy_ddio_ras_n[1] ),
	.phy_ddio_ras_n_2(\phy_ddio_ras_n[2] ),
	.phy_ddio_ras_n_3(\phy_ddio_ras_n[3] ),
	.phy_ddio_reset_n_0(\phy_ddio_reset_n[0] ),
	.phy_ddio_reset_n_1(\phy_ddio_reset_n[1] ),
	.phy_ddio_reset_n_2(\phy_ddio_reset_n[2] ),
	.phy_ddio_reset_n_3(\phy_ddio_reset_n[3] ),
	.phy_ddio_we_n_0(\phy_ddio_we_n[0] ),
	.phy_ddio_we_n_1(\phy_ddio_we_n[1] ),
	.phy_ddio_we_n_2(\phy_ddio_we_n[2] ),
	.phy_ddio_we_n_3(\phy_ddio_we_n[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.ddio_phy_dqslogic_rdatavalid({ddio_phy_dqslogic_rdatavalid_unconnected_wire_4,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_acv_ldc_25 memphy_ldc(
	.pll_dqs_clk(afi_clk),
	.pll_hr_clk(afi_clk),
	.afi_clk(ctl_clk),
	.avl_clk(\memphy_ldc|leveled_hr_clocks[0] ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_mem_phy hphy_inst(
	.aficasn(afi_cas_n[0]),
	.afimemclkdisable(afi_mem_clk_disable[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.avlread(gnd),
	.avlresetn(gnd),
	.avlwrite(gnd),
	.globalresetn(gnd),
	.iointcasnaclr(gnd),
	.iointrasnaclr(gnd),
	.iointresetnaclr(gnd),
	.iointwenaclr(gnd),
	.plladdrcmdclk(!ctl_clk),
	.pllaficlk(ctl_clk),
	.pllavlclk(\memphy_ldc|leveled_hr_clocks[0] ),
	.plllocked(gnd),
	.scanen(gnd),
	.softresetn(gnd),
	.afiaddr({afi_addr[19],afi_addr[18],afi_addr[17],afi_addr[16],afi_addr[15],afi_addr[14],afi_addr[13],afi_addr[12],afi_addr[11],afi_addr[10],afi_addr[9],afi_addr[8],afi_addr[7],afi_addr[6],afi_addr[5],afi_addr[4],afi_addr[3],afi_addr[2],afi_addr[1],afi_addr[0]}),
	.afiba({afi_ba[2],afi_ba[1],afi_ba[0]}),
	.aficke({afi_cke[1],afi_cke[0]}),
	.aficsn({afi_cs_n[1],afi_cs_n[0]}),
	.afidm({afi_dm[9],afi_dm[8],afi_dm[7],afi_dm[6],afi_dm[5],afi_dm[4],afi_dm[3],afi_dm[2],afi_dm[1],afi_dm[0]}),
	.afidqsburst({afi_dqs_burst[4],afi_dqs_burst[3],afi_dqs_burst[2],afi_dqs_burst[1],afi_dqs_burst[0]}),
	.afiodt({afi_odt[1],afi_odt[0]}),
	.afirdataen({afi_rdata_en[4],afi_rdata_en[3],afi_rdata_en[2],afi_rdata_en[1],afi_rdata_en[0]}),
	.afirdataenfull({afi_rdata_en_full[4],afi_rdata_en_full[3],afi_rdata_en_full[2],afi_rdata_en_full[1],afi_rdata_en_full[0]}),
	.afiwdata({afi_wdata[79],afi_wdata[78],afi_wdata[77],afi_wdata[76],afi_wdata[75],afi_wdata[74],afi_wdata[73],afi_wdata[72],afi_wdata[71],afi_wdata[70],afi_wdata[69],afi_wdata[68],afi_wdata[67],afi_wdata[66],afi_wdata[65],afi_wdata[64],afi_wdata[63],afi_wdata[62],afi_wdata[61],afi_wdata[60],afi_wdata[59],afi_wdata[58],afi_wdata[57],afi_wdata[56],afi_wdata[55],afi_wdata[54],afi_wdata[53],afi_wdata[52],
afi_wdata[51],afi_wdata[50],afi_wdata[49],afi_wdata[48],afi_wdata[47],afi_wdata[46],afi_wdata[45],afi_wdata[44],afi_wdata[43],afi_wdata[42],afi_wdata[41],afi_wdata[40],afi_wdata[39],afi_wdata[38],afi_wdata[37],afi_wdata[36],afi_wdata[35],afi_wdata[34],afi_wdata[33],afi_wdata[32],afi_wdata[31],afi_wdata[30],afi_wdata[29],afi_wdata[28],afi_wdata[27],afi_wdata[26],afi_wdata[25],afi_wdata[24],
afi_wdata[23],afi_wdata[22],afi_wdata[21],afi_wdata[20],afi_wdata[19],afi_wdata[18],afi_wdata[17],afi_wdata[16],afi_wdata[15],afi_wdata[14],afi_wdata[13],afi_wdata[12],afi_wdata[11],afi_wdata[10],afi_wdata[9],afi_wdata[8],afi_wdata[7],afi_wdata[6],afi_wdata[5],afi_wdata[4],afi_wdata[3],afi_wdata[2],afi_wdata[1],afi_wdata[0]}),
	.afiwdatavalid({afi_wdata_valid[4],afi_wdata_valid[3],afi_wdata_valid[2],afi_wdata_valid[1],afi_wdata_valid[0]}),
	.avladdress({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.avlwritedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfgaddlat({gnd,gnd,gnd,cfg_addlat[4],cfg_addlat[3],cfg_addlat[2],cfg_addlat[1],cfg_addlat[0]}),
	.cfgbankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth[2],cfg_bankaddrwidth[1],cfg_bankaddrwidth[0]}),
	.cfgcaswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat[3],cfg_caswrlat[2],cfg_caswrlat[1],cfg_caswrlat[0]}),
	.cfgcoladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth[4],cfg_coladdrwidth[3],cfg_coladdrwidth[2],cfg_coladdrwidth[1],cfg_coladdrwidth[0]}),
	.cfgcsaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth[2],cfg_csaddrwidth[1],cfg_csaddrwidth[0]}),
	.cfgdevicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth[3],cfg_devicewidth[2],cfg_devicewidth[1],cfg_devicewidth[0]}),
	.cfgdramconfig({gnd,gnd,gnd,cfg_dramconfig[20],cfg_dramconfig[19],cfg_dramconfig[18],cfg_dramconfig[17],cfg_dramconfig[16],cfg_dramconfig[15],cfg_dramconfig[14],cfg_dramconfig[13],cfg_dramconfig[12],cfg_dramconfig[11],cfg_dramconfig[10],cfg_dramconfig[9],cfg_dramconfig[8],cfg_dramconfig[7],cfg_dramconfig[6],cfg_dramconfig[5],cfg_dramconfig[4],
cfg_dramconfig[3],cfg_dramconfig[2],cfg_dramconfig[1],cfg_dramconfig[0]}),
	.cfginterfacewidth({cfg_interfacewidth[7],cfg_interfacewidth[6],cfg_interfacewidth[5],cfg_interfacewidth[4],cfg_interfacewidth[3],cfg_interfacewidth[2],cfg_interfacewidth[1],cfg_interfacewidth[0]}),
	.cfgrowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth[4],cfg_rowaddrwidth[3],cfg_rowaddrwidth[2],cfg_rowaddrwidth[1],cfg_rowaddrwidth[0]}),
	.cfgtcl({gnd,gnd,gnd,cfg_tcl[4],cfg_tcl[3],cfg_tcl[2],cfg_tcl[1],cfg_tcl[0]}),
	.cfgtmrd({gnd,gnd,gnd,gnd,cfg_tmrd[3],cfg_tmrd[2],cfg_tmrd[1],cfg_tmrd[0]}),
	.cfgtrefi({gnd,gnd,gnd,cfg_trefi[12],cfg_trefi[11],cfg_trefi[10],cfg_trefi[9],cfg_trefi[8],cfg_trefi[7],cfg_trefi[6],cfg_trefi[5],cfg_trefi[4],cfg_trefi[3],cfg_trefi[2],cfg_trefi[1],cfg_trefi[0]}),
	.cfgtrfc({cfg_trfc[7],cfg_trfc[6],cfg_trfc[5],cfg_trfc[4],cfg_trfc[3],cfg_trfc[2],cfg_trfc[1],cfg_trfc[0]}),
	.cfgtwr({gnd,gnd,gnd,gnd,cfg_twr[3],cfg_twr[2],cfg_twr[1],cfg_twr[0]}),
	.ddiophydqdin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] }),
	.ddiophydqslogicrdatavalid({vcc,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.iointaddraclr(16'b0000000000000000),
	.iointaddrdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointbaaclr(3'b000),
	.iointbadout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointcasndout({gnd,gnd,gnd,gnd}),
	.iointckdout({gnd,gnd,gnd,gnd}),
	.iointckeaclr(2'b00),
	.iointckedout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointckndout({gnd,gnd,gnd,gnd}),
	.iointcsnaclr(2'b00),
	.iointcsndout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdmdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iointdqsbdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsboe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicaclrfifoctrl(5'b00000),
	.iointdqslogicaclrpstamble(5'b00000),
	.iointdqslogicdqsena({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicfiforeset({gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincrdataen({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincwrptr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicoct({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicreadlatency({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointodtaclr(2'b00),
	.iointodtdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointrasndout({gnd,gnd,gnd,gnd}),
	.iointresetndout({gnd,gnd,gnd,gnd}),
	.iointwendout({gnd,gnd,gnd,gnd}),
	.aficalfail(afi_cal_fail),
	.aficalsuccess(afi_cal_success),
	.afirdatavalid(afi_rdata_valid[0]),
	.avlwaitrequest(),
	.ctlresetn(ctl_reset_n),
	.iointaficalfail(),
	.iointaficalsuccess(),
	.phyddiocasnaclr(),
	.phyddiorasnaclr(),
	.phyddioresetnaclr(),
	.phyddiowenaclr(),
	.phyresetn(),
	.afirdata(hphy_inst_AFIRDATA_bus),
	.afirlat(),
	.afiwlat(hphy_inst_AFIWLAT_bus),
	.avlreaddata(),
	.iointafirlat(),
	.iointafiwlat(),
	.iointdqdin(),
	.iointdqslogicrdatavalid(),
	.phyddioaddraclr(),
	.phyddioaddrdout(hphy_inst_PHYDDIOADDRDOUT_bus),
	.phyddiobaaclr(),
	.phyddiobadout(hphy_inst_PHYDDIOBADOUT_bus),
	.phyddiocasndout(hphy_inst_PHYDDIOCASNDOUT_bus),
	.phyddiockdout(hphy_inst_PHYDDIOCKDOUT_bus),
	.phyddiockeaclr(),
	.phyddiockedout(hphy_inst_PHYDDIOCKEDOUT_bus),
	.phyddiockndout(),
	.phyddiocsnaclr(),
	.phyddiocsndout(hphy_inst_PHYDDIOCSNDOUT_bus),
	.phyddiodmdout(hphy_inst_PHYDDIODMDOUT_bus),
	.phyddiodqdout(hphy_inst_PHYDDIODQDOUT_bus),
	.phyddiodqoe(hphy_inst_PHYDDIODQOE_bus),
	.phyddiodqsbdout(),
	.phyddiodqsboe(),
	.phyddiodqsdout(hphy_inst_PHYDDIODQSDOUT_bus),
	.phyddiodqslogicaclrfifoctrl(hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus),
	.phyddiodqslogicaclrpstamble(hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus),
	.phyddiodqslogicdqsena(hphy_inst_PHYDDIODQSLOGICDQSENA_bus),
	.phyddiodqslogicfiforeset(hphy_inst_PHYDDIODQSLOGICFIFORESET_bus),
	.phyddiodqslogicincrdataen(hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus),
	.phyddiodqslogicincwrptr(hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus),
	.phyddiodqslogicoct(hphy_inst_PHYDDIODQSLOGICOCT_bus),
	.phyddiodqslogicreadlatency(hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus),
	.phyddiodqsoe(hphy_inst_PHYDDIODQSOE_bus),
	.phyddioodtaclr(),
	.phyddioodtdout(hphy_inst_PHYDDIOODTDOUT_bus),
	.phyddiorasndout(hphy_inst_PHYDDIORASNDOUT_bus),
	.phyddioresetndout(hphy_inst_PHYDDIORESETNDOUT_bus),
	.phyddiowendout(hphy_inst_PHYDDIOWENDOUT_bus));
defparam hphy_inst.hphy_ac_ddr_disable = "true";
defparam hphy_inst.hphy_atpg_en = "false";
defparam hphy_inst.hphy_csr_pipelineglobalenable = "true";
defparam hphy_inst.hphy_datapath_ac_delay = "one_and_half_cycles";
defparam hphy_inst.hphy_datapath_delay = "one_cycle";
defparam hphy_inst.hphy_reset_delay_en = "false";
defparam hphy_inst.hphy_use_hphy = "true";
defparam hphy_inst.hphy_wrap_back_en = "false";
defparam hphy_inst.m_hphy_ac_rom_content = 1200'b100000011100000000000000000000100000011110000000000000000000010000000010000000010001110001010000000010000000010101110000010000000010010000000000000110010000000010100000001000011000010000000010110000000000000000010000001110000000010000000000010000000010000000010001101001010000000010000000010011101000010000000010100000000000000110010000000010010000001000011000010000000010110000000000000000110000011110000000000000000000111000011110000000000000000000110000011110000000000000000000010000011010000000000000000000010000011010110000000000000000010000001010000000010000000000010000010010000000000000000000011100100110000000000000000000011100100110110000000000000000011100100110000000000000001000011100100110110000000000001000111000111110000000000000000000111100111110000000000000000000111000011110000000000000000000011000000110000000000000000000011000100110000000000000000000010011010110000000000000000000010011010110110000000000000000010011010110000000000000001000010011010110110000000000001000110011011110000000000000000000010000010110000000000000001000010000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam hphy_inst.m_hphy_ac_rom_init_file = "hps_ac_rom.hex";
defparam hphy_inst.m_hphy_inst_rom_content = 2560'b1000000000000000000010000000011010000000000010000001100000000000100000100000000000001000001010000000000010000011000000000000100000111000000000001000000100000000000010000100100000000000100001010000000000001000010110000000000010000110000000000000100001000000000000000000100000000000000010000110100000000000000010001000000000001010011010000000100000000110100000000000000010010000000010000000011010000000000000001001100000000000101001101000000000001000011010000000100000000110100000000000000010110110100000001100110011101000000000001010111010000000100011001110100000000000101110001000000011101100100010000000000010100000100000001010110010001000100000000110100000000000110011100000000000001100110110000000000011100111000000000000000011000000000000100000110011100000001000001100111000000010000011001110000000100000110011100000000000001101000000000000000001101000000000000000011010000000000000000110100000000000000001101000000001100000111010000000011000010000100000000110000100001000000001100001000010000000000010100110100000000000100001101000000010000000011010000000000011001110000000000000110011011000000000001110011100000000000000001100000000000011000011001110000000110000110011100000001100001100111000000011000011001110000000000000110100000000000000000110100000000000000001101000000000000000011010000000000000000110100000000111000011101000000001110001000010000000011100010000100000000111000100001000000000001010011010000000000010000110100000001000000001101000000000000001000101011000000000000110110110001000000001101000000000000001000101101000000000000111111010000000000001111110100000001000011111101000010000001111111010000100000100001110100001000001000011101000010000010000111010000000000100010110100000000000011111101000000000000111111010000000101001111110100010000000011010000000010000001110100010000100000100001000100001000001000010001000010000010000100010000100000011110110100001000001000011101000010000010000111010000100000100001110100000001010011010000000010000001111111010000100000100001110100001000001000011101000010000010000111010000100000100000000100001000001000010001000010000010000100010000100000100001000100000000001000100000000000011000110100000000000100001101000000000001110011010000000100000000110100000000000000000000000000000001000000000000000000010100000000000000000110000000000000010000000000000000000000000000000100000000000100000001000000000001010000010000000000011000000100000001000000000001000000000001001000110000000000010000110100000000000101001101000000010000000011010000000010000001111000010001000000001101000000000000000000000000000;
defparam hphy_inst.m_hphy_inst_rom_init_file = "hps_inst_rom.hex";

endmodule

module Computer_System_hps_sdram_p0_acv_hard_io_pads (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	input_path_gen0read_fifo_out_01,
	input_path_gen0read_fifo_out_11,
	input_path_gen0read_fifo_out_21,
	input_path_gen0read_fifo_out_31,
	input_path_gen1read_fifo_out_01,
	input_path_gen1read_fifo_out_11,
	input_path_gen1read_fifo_out_21,
	input_path_gen1read_fifo_out_31,
	input_path_gen2read_fifo_out_01,
	input_path_gen2read_fifo_out_11,
	input_path_gen2read_fifo_out_21,
	input_path_gen2read_fifo_out_31,
	input_path_gen3read_fifo_out_01,
	input_path_gen3read_fifo_out_11,
	input_path_gen3read_fifo_out_21,
	input_path_gen3read_fifo_out_31,
	input_path_gen4read_fifo_out_01,
	input_path_gen4read_fifo_out_11,
	input_path_gen4read_fifo_out_21,
	input_path_gen4read_fifo_out_31,
	input_path_gen5read_fifo_out_01,
	input_path_gen5read_fifo_out_11,
	input_path_gen5read_fifo_out_21,
	input_path_gen5read_fifo_out_31,
	input_path_gen6read_fifo_out_01,
	input_path_gen6read_fifo_out_11,
	input_path_gen6read_fifo_out_21,
	input_path_gen6read_fifo_out_31,
	input_path_gen7read_fifo_out_01,
	input_path_gen7read_fifo_out_11,
	input_path_gen7read_fifo_out_21,
	input_path_gen7read_fifo_out_31,
	input_path_gen0read_fifo_out_02,
	input_path_gen0read_fifo_out_12,
	input_path_gen0read_fifo_out_22,
	input_path_gen0read_fifo_out_32,
	input_path_gen1read_fifo_out_02,
	input_path_gen1read_fifo_out_12,
	input_path_gen1read_fifo_out_22,
	input_path_gen1read_fifo_out_32,
	input_path_gen2read_fifo_out_02,
	input_path_gen2read_fifo_out_12,
	input_path_gen2read_fifo_out_22,
	input_path_gen2read_fifo_out_32,
	input_path_gen3read_fifo_out_02,
	input_path_gen3read_fifo_out_12,
	input_path_gen3read_fifo_out_22,
	input_path_gen3read_fifo_out_32,
	input_path_gen4read_fifo_out_02,
	input_path_gen4read_fifo_out_12,
	input_path_gen4read_fifo_out_22,
	input_path_gen4read_fifo_out_32,
	input_path_gen5read_fifo_out_02,
	input_path_gen5read_fifo_out_12,
	input_path_gen5read_fifo_out_22,
	input_path_gen5read_fifo_out_32,
	input_path_gen6read_fifo_out_02,
	input_path_gen6read_fifo_out_12,
	input_path_gen6read_fifo_out_22,
	input_path_gen6read_fifo_out_32,
	input_path_gen7read_fifo_out_02,
	input_path_gen7read_fifo_out_12,
	input_path_gen7read_fifo_out_22,
	input_path_gen7read_fifo_out_32,
	input_path_gen0read_fifo_out_03,
	input_path_gen0read_fifo_out_13,
	input_path_gen0read_fifo_out_23,
	input_path_gen0read_fifo_out_33,
	input_path_gen1read_fifo_out_03,
	input_path_gen1read_fifo_out_13,
	input_path_gen1read_fifo_out_23,
	input_path_gen1read_fifo_out_33,
	input_path_gen2read_fifo_out_03,
	input_path_gen2read_fifo_out_13,
	input_path_gen2read_fifo_out_23,
	input_path_gen2read_fifo_out_33,
	input_path_gen3read_fifo_out_03,
	input_path_gen3read_fifo_out_13,
	input_path_gen3read_fifo_out_23,
	input_path_gen3read_fifo_out_33,
	input_path_gen4read_fifo_out_03,
	input_path_gen4read_fifo_out_13,
	input_path_gen4read_fifo_out_23,
	input_path_gen4read_fifo_out_33,
	input_path_gen5read_fifo_out_03,
	input_path_gen5read_fifo_out_13,
	input_path_gen5read_fifo_out_23,
	input_path_gen5read_fifo_out_33,
	input_path_gen6read_fifo_out_03,
	input_path_gen6read_fifo_out_13,
	input_path_gen6read_fifo_out_23,
	input_path_gen6read_fifo_out_33,
	input_path_gen7read_fifo_out_03,
	input_path_gen7read_fifo_out_13,
	input_path_gen7read_fifo_out_23,
	input_path_gen7read_fifo_out_33,
	ddio_phy_dqslogic_rdatavalid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	input_path_gen0read_fifo_out_01;
output 	input_path_gen0read_fifo_out_11;
output 	input_path_gen0read_fifo_out_21;
output 	input_path_gen0read_fifo_out_31;
output 	input_path_gen1read_fifo_out_01;
output 	input_path_gen1read_fifo_out_11;
output 	input_path_gen1read_fifo_out_21;
output 	input_path_gen1read_fifo_out_31;
output 	input_path_gen2read_fifo_out_01;
output 	input_path_gen2read_fifo_out_11;
output 	input_path_gen2read_fifo_out_21;
output 	input_path_gen2read_fifo_out_31;
output 	input_path_gen3read_fifo_out_01;
output 	input_path_gen3read_fifo_out_11;
output 	input_path_gen3read_fifo_out_21;
output 	input_path_gen3read_fifo_out_31;
output 	input_path_gen4read_fifo_out_01;
output 	input_path_gen4read_fifo_out_11;
output 	input_path_gen4read_fifo_out_21;
output 	input_path_gen4read_fifo_out_31;
output 	input_path_gen5read_fifo_out_01;
output 	input_path_gen5read_fifo_out_11;
output 	input_path_gen5read_fifo_out_21;
output 	input_path_gen5read_fifo_out_31;
output 	input_path_gen6read_fifo_out_01;
output 	input_path_gen6read_fifo_out_11;
output 	input_path_gen6read_fifo_out_21;
output 	input_path_gen6read_fifo_out_31;
output 	input_path_gen7read_fifo_out_01;
output 	input_path_gen7read_fifo_out_11;
output 	input_path_gen7read_fifo_out_21;
output 	input_path_gen7read_fifo_out_31;
output 	input_path_gen0read_fifo_out_02;
output 	input_path_gen0read_fifo_out_12;
output 	input_path_gen0read_fifo_out_22;
output 	input_path_gen0read_fifo_out_32;
output 	input_path_gen1read_fifo_out_02;
output 	input_path_gen1read_fifo_out_12;
output 	input_path_gen1read_fifo_out_22;
output 	input_path_gen1read_fifo_out_32;
output 	input_path_gen2read_fifo_out_02;
output 	input_path_gen2read_fifo_out_12;
output 	input_path_gen2read_fifo_out_22;
output 	input_path_gen2read_fifo_out_32;
output 	input_path_gen3read_fifo_out_02;
output 	input_path_gen3read_fifo_out_12;
output 	input_path_gen3read_fifo_out_22;
output 	input_path_gen3read_fifo_out_32;
output 	input_path_gen4read_fifo_out_02;
output 	input_path_gen4read_fifo_out_12;
output 	input_path_gen4read_fifo_out_22;
output 	input_path_gen4read_fifo_out_32;
output 	input_path_gen5read_fifo_out_02;
output 	input_path_gen5read_fifo_out_12;
output 	input_path_gen5read_fifo_out_22;
output 	input_path_gen5read_fifo_out_32;
output 	input_path_gen6read_fifo_out_02;
output 	input_path_gen6read_fifo_out_12;
output 	input_path_gen6read_fifo_out_22;
output 	input_path_gen6read_fifo_out_32;
output 	input_path_gen7read_fifo_out_02;
output 	input_path_gen7read_fifo_out_12;
output 	input_path_gen7read_fifo_out_22;
output 	input_path_gen7read_fifo_out_32;
output 	input_path_gen0read_fifo_out_03;
output 	input_path_gen0read_fifo_out_13;
output 	input_path_gen0read_fifo_out_23;
output 	input_path_gen0read_fifo_out_33;
output 	input_path_gen1read_fifo_out_03;
output 	input_path_gen1read_fifo_out_13;
output 	input_path_gen1read_fifo_out_23;
output 	input_path_gen1read_fifo_out_33;
output 	input_path_gen2read_fifo_out_03;
output 	input_path_gen2read_fifo_out_13;
output 	input_path_gen2read_fifo_out_23;
output 	input_path_gen2read_fifo_out_33;
output 	input_path_gen3read_fifo_out_03;
output 	input_path_gen3read_fifo_out_13;
output 	input_path_gen3read_fifo_out_23;
output 	input_path_gen3read_fifo_out_33;
output 	input_path_gen4read_fifo_out_03;
output 	input_path_gen4read_fifo_out_13;
output 	input_path_gen4read_fifo_out_23;
output 	input_path_gen4read_fifo_out_33;
output 	input_path_gen5read_fifo_out_03;
output 	input_path_gen5read_fifo_out_13;
output 	input_path_gen5read_fifo_out_23;
output 	input_path_gen5read_fifo_out_33;
output 	input_path_gen6read_fifo_out_03;
output 	input_path_gen6read_fifo_out_13;
output 	input_path_gen6read_fifo_out_23;
output 	input_path_gen6read_fifo_out_33;
output 	input_path_gen7read_fifo_out_03;
output 	input_path_gen7read_fifo_out_13;
output 	input_path_gen7read_fifo_out_23;
output 	input_path_gen7read_fifo_out_33;
output 	[4:0] ddio_phy_dqslogic_rdatavalid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_hps_sdram_p0_acv_hard_addr_cmd_pads uaddr_cmd_pads(
	.afi_clk(afi_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(phy_ddio_address_0),
	.phy_ddio_address_1(phy_ddio_address_1),
	.phy_ddio_address_2(phy_ddio_address_2),
	.phy_ddio_address_3(phy_ddio_address_3),
	.phy_ddio_address_4(phy_ddio_address_4),
	.phy_ddio_address_5(phy_ddio_address_5),
	.phy_ddio_address_6(phy_ddio_address_6),
	.phy_ddio_address_7(phy_ddio_address_7),
	.phy_ddio_address_8(phy_ddio_address_8),
	.phy_ddio_address_9(phy_ddio_address_9),
	.phy_ddio_address_10(phy_ddio_address_10),
	.phy_ddio_address_11(phy_ddio_address_11),
	.phy_ddio_address_12(phy_ddio_address_12),
	.phy_ddio_address_13(phy_ddio_address_13),
	.phy_ddio_address_14(phy_ddio_address_14),
	.phy_ddio_address_15(phy_ddio_address_15),
	.phy_ddio_address_16(phy_ddio_address_16),
	.phy_ddio_address_17(phy_ddio_address_17),
	.phy_ddio_address_18(phy_ddio_address_18),
	.phy_ddio_address_19(phy_ddio_address_19),
	.phy_ddio_address_20(phy_ddio_address_20),
	.phy_ddio_address_21(phy_ddio_address_21),
	.phy_ddio_address_22(phy_ddio_address_22),
	.phy_ddio_address_23(phy_ddio_address_23),
	.phy_ddio_address_24(phy_ddio_address_24),
	.phy_ddio_address_25(phy_ddio_address_25),
	.phy_ddio_address_26(phy_ddio_address_26),
	.phy_ddio_address_27(phy_ddio_address_27),
	.phy_ddio_address_28(phy_ddio_address_28),
	.phy_ddio_address_29(phy_ddio_address_29),
	.phy_ddio_address_30(phy_ddio_address_30),
	.phy_ddio_address_31(phy_ddio_address_31),
	.phy_ddio_address_32(phy_ddio_address_32),
	.phy_ddio_address_33(phy_ddio_address_33),
	.phy_ddio_address_34(phy_ddio_address_34),
	.phy_ddio_address_35(phy_ddio_address_35),
	.phy_ddio_address_36(phy_ddio_address_36),
	.phy_ddio_address_37(phy_ddio_address_37),
	.phy_ddio_address_38(phy_ddio_address_38),
	.phy_ddio_address_39(phy_ddio_address_39),
	.phy_ddio_address_40(phy_ddio_address_40),
	.phy_ddio_address_41(phy_ddio_address_41),
	.phy_ddio_address_42(phy_ddio_address_42),
	.phy_ddio_address_43(phy_ddio_address_43),
	.phy_ddio_address_44(phy_ddio_address_44),
	.phy_ddio_address_45(phy_ddio_address_45),
	.phy_ddio_address_46(phy_ddio_address_46),
	.phy_ddio_address_47(phy_ddio_address_47),
	.phy_ddio_address_48(phy_ddio_address_48),
	.phy_ddio_address_49(phy_ddio_address_49),
	.phy_ddio_address_50(phy_ddio_address_50),
	.phy_ddio_address_51(phy_ddio_address_51),
	.phy_ddio_address_52(phy_ddio_address_52),
	.phy_ddio_address_53(phy_ddio_address_53),
	.phy_ddio_address_54(phy_ddio_address_54),
	.phy_ddio_address_55(phy_ddio_address_55),
	.phy_ddio_address_56(phy_ddio_address_56),
	.phy_ddio_address_57(phy_ddio_address_57),
	.phy_ddio_address_58(phy_ddio_address_58),
	.phy_ddio_address_59(phy_ddio_address_59),
	.phy_ddio_bank_0(phy_ddio_bank_0),
	.phy_ddio_bank_1(phy_ddio_bank_1),
	.phy_ddio_bank_2(phy_ddio_bank_2),
	.phy_ddio_bank_3(phy_ddio_bank_3),
	.phy_ddio_bank_4(phy_ddio_bank_4),
	.phy_ddio_bank_5(phy_ddio_bank_5),
	.phy_ddio_bank_6(phy_ddio_bank_6),
	.phy_ddio_bank_7(phy_ddio_bank_7),
	.phy_ddio_bank_8(phy_ddio_bank_8),
	.phy_ddio_bank_9(phy_ddio_bank_9),
	.phy_ddio_bank_10(phy_ddio_bank_10),
	.phy_ddio_bank_11(phy_ddio_bank_11),
	.phy_ddio_cas_n_0(phy_ddio_cas_n_0),
	.phy_ddio_cas_n_1(phy_ddio_cas_n_1),
	.phy_ddio_cas_n_2(phy_ddio_cas_n_2),
	.phy_ddio_cas_n_3(phy_ddio_cas_n_3),
	.phy_ddio_ck_0(phy_ddio_ck_0),
	.phy_ddio_ck_1(phy_ddio_ck_1),
	.phy_ddio_cke_0(phy_ddio_cke_0),
	.phy_ddio_cke_1(phy_ddio_cke_1),
	.phy_ddio_cke_2(phy_ddio_cke_2),
	.phy_ddio_cke_3(phy_ddio_cke_3),
	.phy_ddio_cs_n_0(phy_ddio_cs_n_0),
	.phy_ddio_cs_n_1(phy_ddio_cs_n_1),
	.phy_ddio_cs_n_2(phy_ddio_cs_n_2),
	.phy_ddio_cs_n_3(phy_ddio_cs_n_3),
	.phy_ddio_odt_0(phy_ddio_odt_0),
	.phy_ddio_odt_1(phy_ddio_odt_1),
	.phy_ddio_odt_2(phy_ddio_odt_2),
	.phy_ddio_odt_3(phy_ddio_odt_3),
	.phy_ddio_ras_n_0(phy_ddio_ras_n_0),
	.phy_ddio_ras_n_1(phy_ddio_ras_n_1),
	.phy_ddio_ras_n_2(phy_ddio_ras_n_2),
	.phy_ddio_ras_n_3(phy_ddio_ras_n_3),
	.phy_ddio_reset_n_0(phy_ddio_reset_n_0),
	.phy_ddio_reset_n_1(phy_ddio_reset_n_1),
	.phy_ddio_reset_n_2(phy_ddio_reset_n_2),
	.phy_ddio_reset_n_3(phy_ddio_reset_n_3),
	.phy_ddio_we_n_0(phy_ddio_we_n_0),
	.phy_ddio_we_n_1(phy_ddio_we_n_1),
	.phy_ddio_we_n_2(phy_ddio_we_n_2),
	.phy_ddio_we_n_3(phy_ddio_we_n_3),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6));

Computer_System_hps_sdram_p0_altdqdqs_1 \dq_ddio[1].ubidir_dq_dqs (
	.dqsin(dqsin2),
	.pad_gen0raw_input(pad_gen0raw_input2),
	.pad_gen1raw_input(pad_gen1raw_input2),
	.pad_gen2raw_input(pad_gen2raw_input2),
	.pad_gen3raw_input(pad_gen3raw_input2),
	.pad_gen4raw_input(pad_gen4raw_input2),
	.pad_gen5raw_input(pad_gen5raw_input2),
	.pad_gen6raw_input(pad_gen6raw_input2),
	.pad_gen7raw_input(pad_gen7raw_input2),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out2),
	.phy_ddio_dmdout_4(phy_ddio_dmdout_4),
	.phy_ddio_dmdout_5(phy_ddio_dmdout_5),
	.phy_ddio_dmdout_6(phy_ddio_dmdout_6),
	.phy_ddio_dmdout_7(phy_ddio_dmdout_7),
	.phy_ddio_dqdout_36(phy_ddio_dqdout_36),
	.phy_ddio_dqdout_37(phy_ddio_dqdout_37),
	.phy_ddio_dqdout_38(phy_ddio_dqdout_38),
	.phy_ddio_dqdout_39(phy_ddio_dqdout_39),
	.phy_ddio_dqdout_40(phy_ddio_dqdout_40),
	.phy_ddio_dqdout_41(phy_ddio_dqdout_41),
	.phy_ddio_dqdout_42(phy_ddio_dqdout_42),
	.phy_ddio_dqdout_43(phy_ddio_dqdout_43),
	.phy_ddio_dqdout_44(phy_ddio_dqdout_44),
	.phy_ddio_dqdout_45(phy_ddio_dqdout_45),
	.phy_ddio_dqdout_46(phy_ddio_dqdout_46),
	.phy_ddio_dqdout_47(phy_ddio_dqdout_47),
	.phy_ddio_dqdout_48(phy_ddio_dqdout_48),
	.phy_ddio_dqdout_49(phy_ddio_dqdout_49),
	.phy_ddio_dqdout_50(phy_ddio_dqdout_50),
	.phy_ddio_dqdout_51(phy_ddio_dqdout_51),
	.phy_ddio_dqdout_52(phy_ddio_dqdout_52),
	.phy_ddio_dqdout_53(phy_ddio_dqdout_53),
	.phy_ddio_dqdout_54(phy_ddio_dqdout_54),
	.phy_ddio_dqdout_55(phy_ddio_dqdout_55),
	.phy_ddio_dqdout_56(phy_ddio_dqdout_56),
	.phy_ddio_dqdout_57(phy_ddio_dqdout_57),
	.phy_ddio_dqdout_58(phy_ddio_dqdout_58),
	.phy_ddio_dqdout_59(phy_ddio_dqdout_59),
	.phy_ddio_dqdout_60(phy_ddio_dqdout_60),
	.phy_ddio_dqdout_61(phy_ddio_dqdout_61),
	.phy_ddio_dqdout_62(phy_ddio_dqdout_62),
	.phy_ddio_dqdout_63(phy_ddio_dqdout_63),
	.phy_ddio_dqdout_64(phy_ddio_dqdout_64),
	.phy_ddio_dqdout_65(phy_ddio_dqdout_65),
	.phy_ddio_dqdout_66(phy_ddio_dqdout_66),
	.phy_ddio_dqdout_67(phy_ddio_dqdout_67),
	.phy_ddio_dqoe_18(phy_ddio_dqoe_18),
	.phy_ddio_dqoe_19(phy_ddio_dqoe_19),
	.phy_ddio_dqoe_20(phy_ddio_dqoe_20),
	.phy_ddio_dqoe_21(phy_ddio_dqoe_21),
	.phy_ddio_dqoe_22(phy_ddio_dqoe_22),
	.phy_ddio_dqoe_23(phy_ddio_dqoe_23),
	.phy_ddio_dqoe_24(phy_ddio_dqoe_24),
	.phy_ddio_dqoe_25(phy_ddio_dqoe_25),
	.phy_ddio_dqoe_26(phy_ddio_dqoe_26),
	.phy_ddio_dqoe_27(phy_ddio_dqoe_27),
	.phy_ddio_dqoe_28(phy_ddio_dqoe_28),
	.phy_ddio_dqoe_29(phy_ddio_dqoe_29),
	.phy_ddio_dqoe_30(phy_ddio_dqoe_30),
	.phy_ddio_dqoe_31(phy_ddio_dqoe_31),
	.phy_ddio_dqoe_32(phy_ddio_dqoe_32),
	.phy_ddio_dqoe_33(phy_ddio_dqoe_33),
	.phy_ddio_dqs_dout_4(phy_ddio_dqs_dout_4),
	.phy_ddio_dqs_dout_5(phy_ddio_dqs_dout_5),
	.phy_ddio_dqs_dout_6(phy_ddio_dqs_dout_6),
	.phy_ddio_dqs_dout_7(phy_ddio_dqs_dout_7),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.phy_ddio_dqslogic_aclr_pstamble_1(phy_ddio_dqslogic_aclr_pstamble_1),
	.phy_ddio_dqslogic_dqsena_2(phy_ddio_dqslogic_dqsena_2),
	.phy_ddio_dqslogic_dqsena_3(phy_ddio_dqslogic_dqsena_3),
	.phy_ddio_dqslogic_fiforeset_1(phy_ddio_dqslogic_fiforeset_1),
	.phy_ddio_dqslogic_incrdataen_2(phy_ddio_dqslogic_incrdataen_2),
	.phy_ddio_dqslogic_incrdataen_3(phy_ddio_dqslogic_incrdataen_3),
	.phy_ddio_dqslogic_incwrptr_2(phy_ddio_dqslogic_incwrptr_2),
	.phy_ddio_dqslogic_incwrptr_3(phy_ddio_dqslogic_incwrptr_3),
	.phy_ddio_dqslogic_oct_2(phy_ddio_dqslogic_oct_2),
	.phy_ddio_dqslogic_oct_3(phy_ddio_dqslogic_oct_3),
	.phy_ddio_dqslogic_readlatency_5(phy_ddio_dqslogic_readlatency_5),
	.phy_ddio_dqslogic_readlatency_6(phy_ddio_dqslogic_readlatency_6),
	.phy_ddio_dqslogic_readlatency_7(phy_ddio_dqslogic_readlatency_7),
	.phy_ddio_dqslogic_readlatency_8(phy_ddio_dqslogic_readlatency_8),
	.phy_ddio_dqslogic_readlatency_9(phy_ddio_dqslogic_readlatency_9),
	.phy_ddio_dqs_oe_2(phy_ddio_dqs_oe_2),
	.phy_ddio_dqs_oe_3(phy_ddio_dqs_oe_3),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_11),
	.delayed_oct(delayed_oct1),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_11),
	.os(os1),
	.os_bar(os_bar1),
	.diff_oe(diff_oe1),
	.diff_oe_bar(diff_oe_bar1),
	.diff_dtc(diff_dtc1),
	.diff_dtc_bar(diff_dtc_bar1),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_01),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_11),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_21),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_31),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_01),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_11),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_21),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_31),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_01),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_11),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_21),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_31),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_01),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_11),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_21),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_31),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_01),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_11),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_21),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_31),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_01),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_11),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_21),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_31),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_01),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_11),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_21),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_31),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_01),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_11),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_21),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_31),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[1]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_altdqdqs \dq_ddio[0].ubidir_dq_dqs (
	.dqsin(dqsin3),
	.pad_gen0raw_input(pad_gen0raw_input3),
	.pad_gen1raw_input(pad_gen1raw_input3),
	.pad_gen2raw_input(pad_gen2raw_input3),
	.pad_gen3raw_input(pad_gen3raw_input3),
	.pad_gen4raw_input(pad_gen4raw_input3),
	.pad_gen5raw_input(pad_gen5raw_input3),
	.pad_gen6raw_input(pad_gen6raw_input3),
	.pad_gen7raw_input(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out3),
	.phy_ddio_dmdout_0(phy_ddio_dmdout_0),
	.phy_ddio_dmdout_1(phy_ddio_dmdout_1),
	.phy_ddio_dmdout_2(phy_ddio_dmdout_2),
	.phy_ddio_dmdout_3(phy_ddio_dmdout_3),
	.phy_ddio_dqdout_0(phy_ddio_dqdout_0),
	.phy_ddio_dqdout_1(phy_ddio_dqdout_1),
	.phy_ddio_dqdout_2(phy_ddio_dqdout_2),
	.phy_ddio_dqdout_3(phy_ddio_dqdout_3),
	.phy_ddio_dqdout_4(phy_ddio_dqdout_4),
	.phy_ddio_dqdout_5(phy_ddio_dqdout_5),
	.phy_ddio_dqdout_6(phy_ddio_dqdout_6),
	.phy_ddio_dqdout_7(phy_ddio_dqdout_7),
	.phy_ddio_dqdout_8(phy_ddio_dqdout_8),
	.phy_ddio_dqdout_9(phy_ddio_dqdout_9),
	.phy_ddio_dqdout_10(phy_ddio_dqdout_10),
	.phy_ddio_dqdout_11(phy_ddio_dqdout_11),
	.phy_ddio_dqdout_12(phy_ddio_dqdout_12),
	.phy_ddio_dqdout_13(phy_ddio_dqdout_13),
	.phy_ddio_dqdout_14(phy_ddio_dqdout_14),
	.phy_ddio_dqdout_15(phy_ddio_dqdout_15),
	.phy_ddio_dqdout_16(phy_ddio_dqdout_16),
	.phy_ddio_dqdout_17(phy_ddio_dqdout_17),
	.phy_ddio_dqdout_18(phy_ddio_dqdout_18),
	.phy_ddio_dqdout_19(phy_ddio_dqdout_19),
	.phy_ddio_dqdout_20(phy_ddio_dqdout_20),
	.phy_ddio_dqdout_21(phy_ddio_dqdout_21),
	.phy_ddio_dqdout_22(phy_ddio_dqdout_22),
	.phy_ddio_dqdout_23(phy_ddio_dqdout_23),
	.phy_ddio_dqdout_24(phy_ddio_dqdout_24),
	.phy_ddio_dqdout_25(phy_ddio_dqdout_25),
	.phy_ddio_dqdout_26(phy_ddio_dqdout_26),
	.phy_ddio_dqdout_27(phy_ddio_dqdout_27),
	.phy_ddio_dqdout_28(phy_ddio_dqdout_28),
	.phy_ddio_dqdout_29(phy_ddio_dqdout_29),
	.phy_ddio_dqdout_30(phy_ddio_dqdout_30),
	.phy_ddio_dqdout_31(phy_ddio_dqdout_31),
	.phy_ddio_dqoe_0(phy_ddio_dqoe_0),
	.phy_ddio_dqoe_1(phy_ddio_dqoe_1),
	.phy_ddio_dqoe_2(phy_ddio_dqoe_2),
	.phy_ddio_dqoe_3(phy_ddio_dqoe_3),
	.phy_ddio_dqoe_4(phy_ddio_dqoe_4),
	.phy_ddio_dqoe_5(phy_ddio_dqoe_5),
	.phy_ddio_dqoe_6(phy_ddio_dqoe_6),
	.phy_ddio_dqoe_7(phy_ddio_dqoe_7),
	.phy_ddio_dqoe_8(phy_ddio_dqoe_8),
	.phy_ddio_dqoe_9(phy_ddio_dqoe_9),
	.phy_ddio_dqoe_10(phy_ddio_dqoe_10),
	.phy_ddio_dqoe_11(phy_ddio_dqoe_11),
	.phy_ddio_dqoe_12(phy_ddio_dqoe_12),
	.phy_ddio_dqoe_13(phy_ddio_dqoe_13),
	.phy_ddio_dqoe_14(phy_ddio_dqoe_14),
	.phy_ddio_dqoe_15(phy_ddio_dqoe_15),
	.phy_ddio_dqs_dout_0(phy_ddio_dqs_dout_0),
	.phy_ddio_dqs_dout_1(phy_ddio_dqs_dout_1),
	.phy_ddio_dqs_dout_2(phy_ddio_dqs_dout_2),
	.phy_ddio_dqs_dout_3(phy_ddio_dqs_dout_3),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.phy_ddio_dqslogic_aclr_pstamble_0(phy_ddio_dqslogic_aclr_pstamble_0),
	.phy_ddio_dqslogic_dqsena_0(phy_ddio_dqslogic_dqsena_0),
	.phy_ddio_dqslogic_dqsena_1(phy_ddio_dqslogic_dqsena_1),
	.phy_ddio_dqslogic_fiforeset_0(phy_ddio_dqslogic_fiforeset_0),
	.phy_ddio_dqslogic_incrdataen_0(phy_ddio_dqslogic_incrdataen_0),
	.phy_ddio_dqslogic_incrdataen_1(phy_ddio_dqslogic_incrdataen_1),
	.phy_ddio_dqslogic_incwrptr_0(phy_ddio_dqslogic_incwrptr_0),
	.phy_ddio_dqslogic_incwrptr_1(phy_ddio_dqslogic_incwrptr_1),
	.phy_ddio_dqslogic_oct_0(phy_ddio_dqslogic_oct_0),
	.phy_ddio_dqslogic_oct_1(phy_ddio_dqslogic_oct_1),
	.phy_ddio_dqslogic_readlatency_0(phy_ddio_dqslogic_readlatency_0),
	.phy_ddio_dqslogic_readlatency_1(phy_ddio_dqslogic_readlatency_1),
	.phy_ddio_dqslogic_readlatency_2(phy_ddio_dqslogic_readlatency_2),
	.phy_ddio_dqslogic_readlatency_3(phy_ddio_dqslogic_readlatency_3),
	.phy_ddio_dqslogic_readlatency_4(phy_ddio_dqslogic_readlatency_4),
	.phy_ddio_dqs_oe_0(phy_ddio_dqs_oe_0),
	.phy_ddio_dqs_oe_1(phy_ddio_dqs_oe_1),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_0),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_1),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_2),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_3),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_0),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_1),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_2),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_3),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_0),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_1),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_2),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_3),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_0),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_1),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_2),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_3),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_0),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_1),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_2),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_3),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_0),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_1),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_2),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_3),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_0),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_1),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_2),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_3),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_0),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_1),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_2),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_3),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[0]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_altdqdqs_3 \dq_ddio[3].ubidir_dq_dqs (
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.phy_ddio_dmdout_12(phy_ddio_dmdout_12),
	.phy_ddio_dmdout_13(phy_ddio_dmdout_13),
	.phy_ddio_dmdout_14(phy_ddio_dmdout_14),
	.phy_ddio_dmdout_15(phy_ddio_dmdout_15),
	.phy_ddio_dqdout_108(phy_ddio_dqdout_108),
	.phy_ddio_dqdout_109(phy_ddio_dqdout_109),
	.phy_ddio_dqdout_110(phy_ddio_dqdout_110),
	.phy_ddio_dqdout_111(phy_ddio_dqdout_111),
	.phy_ddio_dqdout_112(phy_ddio_dqdout_112),
	.phy_ddio_dqdout_113(phy_ddio_dqdout_113),
	.phy_ddio_dqdout_114(phy_ddio_dqdout_114),
	.phy_ddio_dqdout_115(phy_ddio_dqdout_115),
	.phy_ddio_dqdout_116(phy_ddio_dqdout_116),
	.phy_ddio_dqdout_117(phy_ddio_dqdout_117),
	.phy_ddio_dqdout_118(phy_ddio_dqdout_118),
	.phy_ddio_dqdout_119(phy_ddio_dqdout_119),
	.phy_ddio_dqdout_120(phy_ddio_dqdout_120),
	.phy_ddio_dqdout_121(phy_ddio_dqdout_121),
	.phy_ddio_dqdout_122(phy_ddio_dqdout_122),
	.phy_ddio_dqdout_123(phy_ddio_dqdout_123),
	.phy_ddio_dqdout_124(phy_ddio_dqdout_124),
	.phy_ddio_dqdout_125(phy_ddio_dqdout_125),
	.phy_ddio_dqdout_126(phy_ddio_dqdout_126),
	.phy_ddio_dqdout_127(phy_ddio_dqdout_127),
	.phy_ddio_dqdout_128(phy_ddio_dqdout_128),
	.phy_ddio_dqdout_129(phy_ddio_dqdout_129),
	.phy_ddio_dqdout_130(phy_ddio_dqdout_130),
	.phy_ddio_dqdout_131(phy_ddio_dqdout_131),
	.phy_ddio_dqdout_132(phy_ddio_dqdout_132),
	.phy_ddio_dqdout_133(phy_ddio_dqdout_133),
	.phy_ddio_dqdout_134(phy_ddio_dqdout_134),
	.phy_ddio_dqdout_135(phy_ddio_dqdout_135),
	.phy_ddio_dqdout_136(phy_ddio_dqdout_136),
	.phy_ddio_dqdout_137(phy_ddio_dqdout_137),
	.phy_ddio_dqdout_138(phy_ddio_dqdout_138),
	.phy_ddio_dqdout_139(phy_ddio_dqdout_139),
	.phy_ddio_dqoe_54(phy_ddio_dqoe_54),
	.phy_ddio_dqoe_55(phy_ddio_dqoe_55),
	.phy_ddio_dqoe_56(phy_ddio_dqoe_56),
	.phy_ddio_dqoe_57(phy_ddio_dqoe_57),
	.phy_ddio_dqoe_58(phy_ddio_dqoe_58),
	.phy_ddio_dqoe_59(phy_ddio_dqoe_59),
	.phy_ddio_dqoe_60(phy_ddio_dqoe_60),
	.phy_ddio_dqoe_61(phy_ddio_dqoe_61),
	.phy_ddio_dqoe_62(phy_ddio_dqoe_62),
	.phy_ddio_dqoe_63(phy_ddio_dqoe_63),
	.phy_ddio_dqoe_64(phy_ddio_dqoe_64),
	.phy_ddio_dqoe_65(phy_ddio_dqoe_65),
	.phy_ddio_dqoe_66(phy_ddio_dqoe_66),
	.phy_ddio_dqoe_67(phy_ddio_dqoe_67),
	.phy_ddio_dqoe_68(phy_ddio_dqoe_68),
	.phy_ddio_dqoe_69(phy_ddio_dqoe_69),
	.phy_ddio_dqs_dout_12(phy_ddio_dqs_dout_12),
	.phy_ddio_dqs_dout_13(phy_ddio_dqs_dout_13),
	.phy_ddio_dqs_dout_14(phy_ddio_dqs_dout_14),
	.phy_ddio_dqs_dout_15(phy_ddio_dqs_dout_15),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.phy_ddio_dqslogic_aclr_pstamble_3(phy_ddio_dqslogic_aclr_pstamble_3),
	.phy_ddio_dqslogic_dqsena_6(phy_ddio_dqslogic_dqsena_6),
	.phy_ddio_dqslogic_dqsena_7(phy_ddio_dqslogic_dqsena_7),
	.phy_ddio_dqslogic_fiforeset_3(phy_ddio_dqslogic_fiforeset_3),
	.phy_ddio_dqslogic_incrdataen_6(phy_ddio_dqslogic_incrdataen_6),
	.phy_ddio_dqslogic_incrdataen_7(phy_ddio_dqslogic_incrdataen_7),
	.phy_ddio_dqslogic_incwrptr_6(phy_ddio_dqslogic_incwrptr_6),
	.phy_ddio_dqslogic_incwrptr_7(phy_ddio_dqslogic_incwrptr_7),
	.phy_ddio_dqslogic_oct_6(phy_ddio_dqslogic_oct_6),
	.phy_ddio_dqslogic_oct_7(phy_ddio_dqslogic_oct_7),
	.phy_ddio_dqslogic_readlatency_15(phy_ddio_dqslogic_readlatency_15),
	.phy_ddio_dqslogic_readlatency_16(phy_ddio_dqslogic_readlatency_16),
	.phy_ddio_dqslogic_readlatency_17(phy_ddio_dqslogic_readlatency_17),
	.phy_ddio_dqslogic_readlatency_18(phy_ddio_dqslogic_readlatency_18),
	.phy_ddio_dqslogic_readlatency_19(phy_ddio_dqslogic_readlatency_19),
	.phy_ddio_dqs_oe_6(phy_ddio_dqs_oe_6),
	.phy_ddio_dqs_oe_7(phy_ddio_dqs_oe_7),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_13),
	.delayed_oct(delayed_oct3),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_13),
	.os(os3),
	.os_bar(os_bar3),
	.diff_oe(diff_oe3),
	.diff_oe_bar(diff_oe_bar3),
	.diff_dtc(diff_dtc3),
	.diff_dtc_bar(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_03),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_13),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_23),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_33),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_03),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_13),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_23),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_33),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_03),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_13),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_23),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_33),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_03),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_13),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_23),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_33),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_03),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_13),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_23),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_33),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_03),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_13),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_23),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_33),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_03),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_13),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_23),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_33),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_03),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_13),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_23),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_33),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[3]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_altdqdqs_2 \dq_ddio[2].ubidir_dq_dqs (
	.dqsin(dqsin1),
	.pad_gen0raw_input(pad_gen0raw_input1),
	.pad_gen1raw_input(pad_gen1raw_input1),
	.pad_gen2raw_input(pad_gen2raw_input1),
	.pad_gen3raw_input(pad_gen3raw_input1),
	.pad_gen4raw_input(pad_gen4raw_input1),
	.pad_gen5raw_input(pad_gen5raw_input1),
	.pad_gen6raw_input(pad_gen6raw_input1),
	.pad_gen7raw_input(pad_gen7raw_input1),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out1),
	.phy_ddio_dmdout_8(phy_ddio_dmdout_8),
	.phy_ddio_dmdout_9(phy_ddio_dmdout_9),
	.phy_ddio_dmdout_10(phy_ddio_dmdout_10),
	.phy_ddio_dmdout_11(phy_ddio_dmdout_11),
	.phy_ddio_dqdout_72(phy_ddio_dqdout_72),
	.phy_ddio_dqdout_73(phy_ddio_dqdout_73),
	.phy_ddio_dqdout_74(phy_ddio_dqdout_74),
	.phy_ddio_dqdout_75(phy_ddio_dqdout_75),
	.phy_ddio_dqdout_76(phy_ddio_dqdout_76),
	.phy_ddio_dqdout_77(phy_ddio_dqdout_77),
	.phy_ddio_dqdout_78(phy_ddio_dqdout_78),
	.phy_ddio_dqdout_79(phy_ddio_dqdout_79),
	.phy_ddio_dqdout_80(phy_ddio_dqdout_80),
	.phy_ddio_dqdout_81(phy_ddio_dqdout_81),
	.phy_ddio_dqdout_82(phy_ddio_dqdout_82),
	.phy_ddio_dqdout_83(phy_ddio_dqdout_83),
	.phy_ddio_dqdout_84(phy_ddio_dqdout_84),
	.phy_ddio_dqdout_85(phy_ddio_dqdout_85),
	.phy_ddio_dqdout_86(phy_ddio_dqdout_86),
	.phy_ddio_dqdout_87(phy_ddio_dqdout_87),
	.phy_ddio_dqdout_88(phy_ddio_dqdout_88),
	.phy_ddio_dqdout_89(phy_ddio_dqdout_89),
	.phy_ddio_dqdout_90(phy_ddio_dqdout_90),
	.phy_ddio_dqdout_91(phy_ddio_dqdout_91),
	.phy_ddio_dqdout_92(phy_ddio_dqdout_92),
	.phy_ddio_dqdout_93(phy_ddio_dqdout_93),
	.phy_ddio_dqdout_94(phy_ddio_dqdout_94),
	.phy_ddio_dqdout_95(phy_ddio_dqdout_95),
	.phy_ddio_dqdout_96(phy_ddio_dqdout_96),
	.phy_ddio_dqdout_97(phy_ddio_dqdout_97),
	.phy_ddio_dqdout_98(phy_ddio_dqdout_98),
	.phy_ddio_dqdout_99(phy_ddio_dqdout_99),
	.phy_ddio_dqdout_100(phy_ddio_dqdout_100),
	.phy_ddio_dqdout_101(phy_ddio_dqdout_101),
	.phy_ddio_dqdout_102(phy_ddio_dqdout_102),
	.phy_ddio_dqdout_103(phy_ddio_dqdout_103),
	.phy_ddio_dqoe_36(phy_ddio_dqoe_36),
	.phy_ddio_dqoe_37(phy_ddio_dqoe_37),
	.phy_ddio_dqoe_38(phy_ddio_dqoe_38),
	.phy_ddio_dqoe_39(phy_ddio_dqoe_39),
	.phy_ddio_dqoe_40(phy_ddio_dqoe_40),
	.phy_ddio_dqoe_41(phy_ddio_dqoe_41),
	.phy_ddio_dqoe_42(phy_ddio_dqoe_42),
	.phy_ddio_dqoe_43(phy_ddio_dqoe_43),
	.phy_ddio_dqoe_44(phy_ddio_dqoe_44),
	.phy_ddio_dqoe_45(phy_ddio_dqoe_45),
	.phy_ddio_dqoe_46(phy_ddio_dqoe_46),
	.phy_ddio_dqoe_47(phy_ddio_dqoe_47),
	.phy_ddio_dqoe_48(phy_ddio_dqoe_48),
	.phy_ddio_dqoe_49(phy_ddio_dqoe_49),
	.phy_ddio_dqoe_50(phy_ddio_dqoe_50),
	.phy_ddio_dqoe_51(phy_ddio_dqoe_51),
	.phy_ddio_dqs_dout_8(phy_ddio_dqs_dout_8),
	.phy_ddio_dqs_dout_9(phy_ddio_dqs_dout_9),
	.phy_ddio_dqs_dout_10(phy_ddio_dqs_dout_10),
	.phy_ddio_dqs_dout_11(phy_ddio_dqs_dout_11),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.phy_ddio_dqslogic_aclr_pstamble_2(phy_ddio_dqslogic_aclr_pstamble_2),
	.phy_ddio_dqslogic_dqsena_4(phy_ddio_dqslogic_dqsena_4),
	.phy_ddio_dqslogic_dqsena_5(phy_ddio_dqslogic_dqsena_5),
	.phy_ddio_dqslogic_fiforeset_2(phy_ddio_dqslogic_fiforeset_2),
	.phy_ddio_dqslogic_incrdataen_4(phy_ddio_dqslogic_incrdataen_4),
	.phy_ddio_dqslogic_incrdataen_5(phy_ddio_dqslogic_incrdataen_5),
	.phy_ddio_dqslogic_incwrptr_4(phy_ddio_dqslogic_incwrptr_4),
	.phy_ddio_dqslogic_incwrptr_5(phy_ddio_dqslogic_incwrptr_5),
	.phy_ddio_dqslogic_oct_4(phy_ddio_dqslogic_oct_4),
	.phy_ddio_dqslogic_oct_5(phy_ddio_dqslogic_oct_5),
	.phy_ddio_dqslogic_readlatency_10(phy_ddio_dqslogic_readlatency_10),
	.phy_ddio_dqslogic_readlatency_11(phy_ddio_dqslogic_readlatency_11),
	.phy_ddio_dqslogic_readlatency_12(phy_ddio_dqslogic_readlatency_12),
	.phy_ddio_dqslogic_readlatency_13(phy_ddio_dqslogic_readlatency_13),
	.phy_ddio_dqslogic_readlatency_14(phy_ddio_dqslogic_readlatency_14),
	.phy_ddio_dqs_oe_4(phy_ddio_dqs_oe_4),
	.phy_ddio_dqs_oe_5(phy_ddio_dqs_oe_5),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_12),
	.delayed_oct(delayed_oct2),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_12),
	.os(os2),
	.os_bar(os_bar2),
	.diff_oe(diff_oe2),
	.diff_oe_bar(diff_oe_bar2),
	.diff_dtc(diff_dtc2),
	.diff_dtc_bar(diff_dtc_bar2),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_02),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_12),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_22),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_32),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_02),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_12),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_22),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_32),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_02),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_12),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_22),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_32),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_02),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_12),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_22),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_32),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_02),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_12),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_22),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_32),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_02),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_12),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_22),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_32),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_02),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_12),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_22),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_32),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_02),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_12),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_22),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_32),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[2]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module Computer_System_hps_sdram_p0_acv_hard_addr_cmd_pads (
	afi_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6)/* synthesis synthesis_greybox=0 */;
input 	afi_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_gen[0].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[1].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[2].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[3].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[4].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[5].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[6].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[7].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[8].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[9].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[10].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[11].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[12].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[13].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[14].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[15].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[16].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[17].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[19].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[18].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[21].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[22].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[23].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[24].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[20].acv_ac_ldc|adc_clk_cps ;
wire \clock_gen[0].umem_ck_pad|auto_generated|dataout[0] ;
wire \mem_ck_source[0] ;
wire \clock_gen[0].leveled_dqs_clocks[0] ;
wire \clock_gen[0].leveled_dqs_clocks[1] ;
wire \clock_gen[0].leveled_dqs_clocks[2] ;
wire \clock_gen[0].leveled_dqs_clocks[3] ;

wire [3:0] \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ;

assign \clock_gen[0].leveled_dqs_clocks[0]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [0];
assign \clock_gen[0].leveled_dqs_clocks[1]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [1];
assign \clock_gen[0].leveled_dqs_clocks[2]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [2];
assign \clock_gen[0].leveled_dqs_clocks[3]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [3];

Computer_System_hps_sdram_p0_acv_ldc_19 \address_gen[4].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[4].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_18 \address_gen[3].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[3].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_17 \address_gen[2].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[2].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_11 \address_gen[1].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[1].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc \address_gen[0].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[0].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_2 \address_gen[11].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[11].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_1 \address_gen[10].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[10].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_24 \address_gen[9].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[9].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_23 \address_gen[8].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[8].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_22 \address_gen[7].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[7].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_21 \address_gen[6].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[6].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_20 \address_gen[5].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[5].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_10 \address_gen[19].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[19].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_9 \address_gen[18].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[18].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_8 \address_gen[17].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[17].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_7 \address_gen[16].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[16].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_6 \address_gen[15].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[15].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_5 \address_gen[14].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[14].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_4 \address_gen[13].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[13].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_3 \address_gen[12].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[12].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_generic_ddio_1 ubank_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14,dataout_unconnected_wire_13,dataout_unconnected_wire_12,dataout_unconnected_wire_11,dataout_unconnected_wire_10,dataout_unconnected_wire_9,dataout_unconnected_wire_8,dataout_unconnected_wire_7,dataout_unconnected_wire_6,
dataout_unconnected_wire_5,dataout_unconnected_wire_4,dataout_unconnected_wire_3,dataout_21,dataout_15,dataout_01}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[17].acv_ac_ldc|adc_clk_cps ,\address_gen[16].acv_ac_ldc|adc_clk_cps ,\address_gen[15].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_bank_11,phy_ddio_bank_10,phy_ddio_bank_9,phy_ddio_bank_8,phy_ddio_bank_7,phy_ddio_bank_6,phy_ddio_bank_5,
phy_ddio_bank_4,phy_ddio_bank_3,phy_ddio_bank_2,phy_ddio_bank_1,phy_ddio_bank_0}));

Computer_System_hps_sdram_p0_generic_ddio uaddress_pad(
	.clk_hr({afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_14,dataout_13,dataout_12,dataout_11,dataout_10,dataout_9,dataout_8,dataout_7,dataout_6,dataout_5,dataout_4,dataout_3,dataout_2,dataout_1,dataout_0}),
	.clk_fr({\address_gen[14].acv_ac_ldc|adc_clk_cps ,\address_gen[13].acv_ac_ldc|adc_clk_cps ,\address_gen[12].acv_ac_ldc|adc_clk_cps ,\address_gen[11].acv_ac_ldc|adc_clk_cps ,\address_gen[10].acv_ac_ldc|adc_clk_cps ,\address_gen[9].acv_ac_ldc|adc_clk_cps ,
\address_gen[8].acv_ac_ldc|adc_clk_cps ,\address_gen[7].acv_ac_ldc|adc_clk_cps ,\address_gen[6].acv_ac_ldc|adc_clk_cps ,\address_gen[5].acv_ac_ldc|adc_clk_cps ,\address_gen[4].acv_ac_ldc|adc_clk_cps ,\address_gen[3].acv_ac_ldc|adc_clk_cps ,
\address_gen[2].acv_ac_ldc|adc_clk_cps ,\address_gen[1].acv_ac_ldc|adc_clk_cps ,\address_gen[0].acv_ac_ldc|adc_clk_cps }),
	.datain({phy_ddio_address_59,phy_ddio_address_58,phy_ddio_address_57,phy_ddio_address_56,phy_ddio_address_55,phy_ddio_address_54,phy_ddio_address_53,phy_ddio_address_52,phy_ddio_address_51,phy_ddio_address_50,phy_ddio_address_49,phy_ddio_address_48,phy_ddio_address_47,
phy_ddio_address_46,phy_ddio_address_45,phy_ddio_address_44,phy_ddio_address_43,phy_ddio_address_42,phy_ddio_address_41,phy_ddio_address_40,phy_ddio_address_39,phy_ddio_address_38,phy_ddio_address_37,phy_ddio_address_36,phy_ddio_address_35,phy_ddio_address_34,
phy_ddio_address_33,phy_ddio_address_32,phy_ddio_address_31,phy_ddio_address_30,phy_ddio_address_29,phy_ddio_address_28,phy_ddio_address_27,phy_ddio_address_26,phy_ddio_address_25,phy_ddio_address_24,phy_ddio_address_23,phy_ddio_address_22,phy_ddio_address_21,
phy_ddio_address_20,phy_ddio_address_19,phy_ddio_address_18,phy_ddio_address_17,phy_ddio_address_16,phy_ddio_address_15,phy_ddio_address_14,phy_ddio_address_13,phy_ddio_address_12,phy_ddio_address_11,phy_ddio_address_10,phy_ddio_address_9,phy_ddio_address_8,
phy_ddio_address_7,phy_ddio_address_6,phy_ddio_address_5,phy_ddio_address_4,phy_ddio_address_3,phy_ddio_address_2,phy_ddio_address_1,phy_ddio_address_0}));

Computer_System_hps_sdram_p0_acv_ldc_16 \address_gen[24].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[24].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_15 \address_gen[23].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[23].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_14 \address_gen[22].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[22].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_13 \address_gen[21].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[21].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_12 \address_gen[20].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[20].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_clock_pair_generator \clock_gen[0].uclk_generator (
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.datain({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }));

Computer_System_altddio_out_1 \clock_gen[0].umem_ck_pad (
	.dataout({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }),
	.datain_h({phy_ddio_ck_0}),
	.datain_l({phy_ddio_ck_1}),
	.outclock(\mem_ck_source[0] ));

Computer_System_hps_sdram_p0_generic_ddio_3 ureset_n_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk}),
	.dataout({dataout_unconnected_wire_14_1,dataout_unconnected_wire_13_1,dataout_unconnected_wire_12_1,dataout_unconnected_wire_11_1,dataout_unconnected_wire_10_1,dataout_unconnected_wire_9_1,dataout_unconnected_wire_8_1,dataout_unconnected_wire_7_1,
dataout_unconnected_wire_6_1,dataout_unconnected_wire_5_1,dataout_unconnected_wire_4_1,dataout_unconnected_wire_3_1,dataout_unconnected_wire_2,dataout_unconnected_wire_1,dataout_03}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[24].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_reset_n_3,phy_ddio_reset_n_2,phy_ddio_reset_n_1,phy_ddio_reset_n_0}));

Computer_System_hps_sdram_p0_generic_ddio_2 ucmd_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_2,dataout_unconnected_wire_13_2,dataout_unconnected_wire_12_2,dataout_unconnected_wire_11_2,dataout_unconnected_wire_10_2,dataout_unconnected_wire_9_2,dataout_unconnected_wire_8_2,dataout_unconnected_wire_7_2,
dataout_unconnected_wire_6_2,dataout_51,dataout_41,dataout_31,dataout_22,dataout_16,dataout_02}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[23].acv_ac_ldc|adc_clk_cps ,\address_gen[22].acv_ac_ldc|adc_clk_cps ,\address_gen[21].acv_ac_ldc|adc_clk_cps ,\address_gen[20].acv_ac_ldc|adc_clk_cps ,\address_gen[19].acv_ac_ldc|adc_clk_cps ,
\address_gen[18].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_we_n_3,phy_ddio_we_n_2,phy_ddio_we_n_1,phy_ddio_we_n_0,phy_ddio_cas_n_3,phy_ddio_cas_n_2,phy_ddio_cas_n_1,phy_ddio_cas_n_0,phy_ddio_ras_n_3,
phy_ddio_ras_n_2,phy_ddio_ras_n_1,phy_ddio_ras_n_0,phy_ddio_odt_3,phy_ddio_odt_2,phy_ddio_odt_1,phy_ddio_odt_0,phy_ddio_cke_3,phy_ddio_cke_2,phy_ddio_cke_1,phy_ddio_cke_0,phy_ddio_cs_n_3,phy_ddio_cs_n_2,phy_ddio_cs_n_1,phy_ddio_cs_n_0}));

cyclonev_clk_phase_select \clock_gen[0].clk_phase_select_dqs (
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\clock_gen[0].leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(\mem_ck_source[0] ));
defparam \clock_gen[0].clk_phase_select_dqs .invert_phase = "false";
defparam \clock_gen[0].clk_phase_select_dqs .phase_setting = 0;
defparam \clock_gen[0].clk_phase_select_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].clk_phase_select_dqs .use_dqs_input = "false";
defparam \clock_gen[0].clk_phase_select_dqs .use_phasectrlin = "false";

cyclonev_leveling_delay_chain \clock_gen[0].leveling_delay_chain_dqs (
	.clkin(afi_clk),
	.delayctrlin({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.clkout(\clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ));
defparam \clock_gen[0].leveling_delay_chain_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_delay_increment = 10;
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_altddio_out_1 (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
inout 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_ddio_out_uqe auto_generated(
	.dataout({dataout[0]}),
	.datain_h({datain_h[0]}),
	.datain_l({datain_l[0]}),
	.outclock(outclock));

endmodule

module Computer_System_ddio_out_uqe (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
output 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "none";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_acv_ldc (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_1 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_2 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_3 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_4 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_5 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_6 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_7 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_8 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_9 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_10 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_11 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_12 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_13 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_14 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_15 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_16 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_17 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_18 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_19 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_20 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_21 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_22 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_23 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_24 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_clock_pair_generator (
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	datain)/* synthesis synthesis_greybox=0 */;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	[0:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(datain[0]),
	.oein(gnd),
	.dtcin(gnd),
	.o(wire_pseudo_diffa_o_0),
	.obar(wire_pseudo_diffa_obar_0),
	.oeout(wire_pseudo_diffa_oeout_0),
	.oebout(wire_pseudo_diffa_oebout_0),
	.dtc(),
	.dtcbar());

endmodule

module Computer_System_hps_sdram_p0_generic_ddio (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[6].fr_data_lo ;
wire \acblock[6].fr_data_hi ;
wire \acblock[7].fr_data_lo ;
wire \acblock[7].fr_data_hi ;
wire \acblock[8].fr_data_lo ;
wire \acblock[8].fr_data_hi ;
wire \acblock[9].fr_data_lo ;
wire \acblock[9].fr_data_hi ;
wire \acblock[10].fr_data_lo ;
wire \acblock[10].fr_data_hi ;
wire \acblock[11].fr_data_lo ;
wire \acblock[11].fr_data_hi ;
wire \acblock[12].fr_data_lo ;
wire \acblock[12].fr_data_hi ;
wire \acblock[13].fr_data_lo ;
wire \acblock[13].fr_data_hi ;
wire \acblock[14].fr_data_lo ;
wire \acblock[14].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].ddio_out (
	.datainlo(\acblock[6].fr_data_lo ),
	.datainhi(\acblock[6].fr_data_hi ),
	.clkhi(clk_fr[6]),
	.clklo(clk_fr[6]),
	.muxsel(clk_fr[6]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[6]),
	.dfflo(),
	.dffhi());
defparam \acblock[6].ddio_out .async_mode = "none";
defparam \acblock[6].ddio_out .half_rate_mode = "false";
defparam \acblock[6].ddio_out .power_up = "low";
defparam \acblock[6].ddio_out .sync_mode = "none";
defparam \acblock[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].ddio_out (
	.datainlo(\acblock[7].fr_data_lo ),
	.datainhi(\acblock[7].fr_data_hi ),
	.clkhi(clk_fr[7]),
	.clklo(clk_fr[7]),
	.muxsel(clk_fr[7]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[7]),
	.dfflo(),
	.dffhi());
defparam \acblock[7].ddio_out .async_mode = "none";
defparam \acblock[7].ddio_out .half_rate_mode = "false";
defparam \acblock[7].ddio_out .power_up = "low";
defparam \acblock[7].ddio_out .sync_mode = "none";
defparam \acblock[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].ddio_out (
	.datainlo(\acblock[8].fr_data_lo ),
	.datainhi(\acblock[8].fr_data_hi ),
	.clkhi(clk_fr[8]),
	.clklo(clk_fr[8]),
	.muxsel(clk_fr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[8]),
	.dfflo(),
	.dffhi());
defparam \acblock[8].ddio_out .async_mode = "none";
defparam \acblock[8].ddio_out .half_rate_mode = "false";
defparam \acblock[8].ddio_out .power_up = "low";
defparam \acblock[8].ddio_out .sync_mode = "none";
defparam \acblock[8].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].ddio_out (
	.datainlo(\acblock[9].fr_data_lo ),
	.datainhi(\acblock[9].fr_data_hi ),
	.clkhi(clk_fr[9]),
	.clklo(clk_fr[9]),
	.muxsel(clk_fr[9]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[9]),
	.dfflo(),
	.dffhi());
defparam \acblock[9].ddio_out .async_mode = "none";
defparam \acblock[9].ddio_out .half_rate_mode = "false";
defparam \acblock[9].ddio_out .power_up = "low";
defparam \acblock[9].ddio_out .sync_mode = "none";
defparam \acblock[9].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].ddio_out (
	.datainlo(\acblock[10].fr_data_lo ),
	.datainhi(\acblock[10].fr_data_hi ),
	.clkhi(clk_fr[10]),
	.clklo(clk_fr[10]),
	.muxsel(clk_fr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[10]),
	.dfflo(),
	.dffhi());
defparam \acblock[10].ddio_out .async_mode = "none";
defparam \acblock[10].ddio_out .half_rate_mode = "false";
defparam \acblock[10].ddio_out .power_up = "low";
defparam \acblock[10].ddio_out .sync_mode = "none";
defparam \acblock[10].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].ddio_out (
	.datainlo(\acblock[11].fr_data_lo ),
	.datainhi(\acblock[11].fr_data_hi ),
	.clkhi(clk_fr[11]),
	.clklo(clk_fr[11]),
	.muxsel(clk_fr[11]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[11]),
	.dfflo(),
	.dffhi());
defparam \acblock[11].ddio_out .async_mode = "none";
defparam \acblock[11].ddio_out .half_rate_mode = "false";
defparam \acblock[11].ddio_out .power_up = "low";
defparam \acblock[11].ddio_out .sync_mode = "none";
defparam \acblock[11].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].ddio_out (
	.datainlo(\acblock[12].fr_data_lo ),
	.datainhi(\acblock[12].fr_data_hi ),
	.clkhi(clk_fr[12]),
	.clklo(clk_fr[12]),
	.muxsel(clk_fr[12]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[12]),
	.dfflo(),
	.dffhi());
defparam \acblock[12].ddio_out .async_mode = "none";
defparam \acblock[12].ddio_out .half_rate_mode = "false";
defparam \acblock[12].ddio_out .power_up = "low";
defparam \acblock[12].ddio_out .sync_mode = "none";
defparam \acblock[12].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].ddio_out (
	.datainlo(\acblock[13].fr_data_lo ),
	.datainhi(\acblock[13].fr_data_hi ),
	.clkhi(clk_fr[13]),
	.clklo(clk_fr[13]),
	.muxsel(clk_fr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[13]),
	.dfflo(),
	.dffhi());
defparam \acblock[13].ddio_out .async_mode = "none";
defparam \acblock[13].ddio_out .half_rate_mode = "false";
defparam \acblock[13].ddio_out .power_up = "low";
defparam \acblock[13].ddio_out .sync_mode = "none";
defparam \acblock[13].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].ddio_out (
	.datainlo(\acblock[14].fr_data_lo ),
	.datainhi(\acblock[14].fr_data_hi ),
	.clkhi(clk_fr[14]),
	.clklo(clk_fr[14]),
	.muxsel(clk_fr[14]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[14]),
	.dfflo(),
	.dffhi());
defparam \acblock[14].ddio_out .async_mode = "none";
defparam \acblock[14].ddio_out .half_rate_mode = "false";
defparam \acblock[14].ddio_out .power_up = "low";
defparam \acblock[14].ddio_out .sync_mode = "none";
defparam \acblock[14].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_lo (
	.datainlo(datain[27]),
	.datainhi(datain[25]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_lo .async_mode = "none";
defparam \acblock[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_lo .power_up = "low";
defparam \acblock[6].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_hi (
	.datainlo(datain[26]),
	.datainhi(datain[24]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_hi .async_mode = "none";
defparam \acblock[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_hi .power_up = "low";
defparam \acblock[6].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_lo (
	.datainlo(datain[31]),
	.datainhi(datain[29]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_lo .async_mode = "none";
defparam \acblock[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_lo .power_up = "low";
defparam \acblock[7].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_hi (
	.datainlo(datain[30]),
	.datainhi(datain[28]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_hi .async_mode = "none";
defparam \acblock[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_hi .power_up = "low";
defparam \acblock[7].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_lo (
	.datainlo(datain[35]),
	.datainhi(datain[33]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_lo .async_mode = "none";
defparam \acblock[8].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_lo .power_up = "low";
defparam \acblock[8].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[8].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_hi (
	.datainlo(datain[34]),
	.datainhi(datain[32]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_hi .async_mode = "none";
defparam \acblock[8].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_hi .power_up = "low";
defparam \acblock[8].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[8].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_lo (
	.datainlo(datain[39]),
	.datainhi(datain[37]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_lo .async_mode = "none";
defparam \acblock[9].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_lo .power_up = "low";
defparam \acblock[9].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[9].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_hi (
	.datainlo(datain[38]),
	.datainhi(datain[36]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_hi .async_mode = "none";
defparam \acblock[9].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_hi .power_up = "low";
defparam \acblock[9].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[9].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_lo (
	.datainlo(datain[43]),
	.datainhi(datain[41]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_lo .async_mode = "none";
defparam \acblock[10].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_lo .power_up = "low";
defparam \acblock[10].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[10].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_hi (
	.datainlo(datain[42]),
	.datainhi(datain[40]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_hi .async_mode = "none";
defparam \acblock[10].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_hi .power_up = "low";
defparam \acblock[10].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[10].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_lo (
	.datainlo(datain[47]),
	.datainhi(datain[45]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_lo .async_mode = "none";
defparam \acblock[11].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_lo .power_up = "low";
defparam \acblock[11].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[11].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_hi (
	.datainlo(datain[46]),
	.datainhi(datain[44]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_hi .async_mode = "none";
defparam \acblock[11].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_hi .power_up = "low";
defparam \acblock[11].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[11].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_lo (
	.datainlo(datain[51]),
	.datainhi(datain[49]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_lo .async_mode = "none";
defparam \acblock[12].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_lo .power_up = "low";
defparam \acblock[12].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[12].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_hi (
	.datainlo(datain[50]),
	.datainhi(datain[48]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_hi .async_mode = "none";
defparam \acblock[12].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_hi .power_up = "low";
defparam \acblock[12].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[12].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_lo (
	.datainlo(datain[55]),
	.datainhi(datain[53]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_lo .async_mode = "none";
defparam \acblock[13].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_lo .power_up = "low";
defparam \acblock[13].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[13].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_hi (
	.datainlo(datain[54]),
	.datainhi(datain[52]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_hi .async_mode = "none";
defparam \acblock[13].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_hi .power_up = "low";
defparam \acblock[13].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[13].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_lo (
	.datainlo(datain[59]),
	.datainhi(datain[57]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_lo .async_mode = "none";
defparam \acblock[14].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_lo .power_up = "low";
defparam \acblock[14].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[14].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_hi (
	.datainlo(datain[58]),
	.datainhi(datain[56]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_hi .async_mode = "none";
defparam \acblock[14].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_hi .power_up = "low";
defparam \acblock[14].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[14].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_generic_ddio_1 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_generic_ddio_2 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_generic_ddio_3 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_3,phy_ddio_dmdout_2,phy_ddio_dmdout_1,phy_ddio_dmdout_0}),
	.write_data_in({phy_ddio_dqdout_31,phy_ddio_dqdout_30,phy_ddio_dqdout_29,phy_ddio_dqdout_28,phy_ddio_dqdout_27,phy_ddio_dqdout_26,phy_ddio_dqdout_25,phy_ddio_dqdout_24,phy_ddio_dqdout_23,phy_ddio_dqdout_22,phy_ddio_dqdout_21,phy_ddio_dqdout_20,phy_ddio_dqdout_19,phy_ddio_dqdout_18,
phy_ddio_dqdout_17,phy_ddio_dqdout_16,phy_ddio_dqdout_15,phy_ddio_dqdout_14,phy_ddio_dqdout_13,phy_ddio_dqdout_12,phy_ddio_dqdout_11,phy_ddio_dqdout_10,phy_ddio_dqdout_9,phy_ddio_dqdout_8,phy_ddio_dqdout_7,phy_ddio_dqdout_6,phy_ddio_dqdout_5,phy_ddio_dqdout_4,
phy_ddio_dqdout_3,phy_ddio_dqdout_2,phy_ddio_dqdout_1,phy_ddio_dqdout_0}),
	.write_oe_in({phy_ddio_dqoe_15,phy_ddio_dqoe_14,phy_ddio_dqoe_13,phy_ddio_dqoe_12,phy_ddio_dqoe_11,phy_ddio_dqoe_10,phy_ddio_dqoe_9,phy_ddio_dqoe_8,phy_ddio_dqoe_7,phy_ddio_dqoe_6,phy_ddio_dqoe_5,phy_ddio_dqoe_4,phy_ddio_dqoe_3,phy_ddio_dqoe_2,phy_ddio_dqoe_1,phy_ddio_dqoe_0}),
	.write_strobe({phy_ddio_dqs_dout_3,phy_ddio_dqs_dout_2,phy_ddio_dqs_dout_1,phy_ddio_dqs_dout_0}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_0),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_0),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_1,phy_ddio_dqslogic_incrdataen_0}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_1,phy_ddio_dqslogic_incwrptr_0}),
	.oct_ena_in({phy_ddio_dqslogic_oct_1,phy_ddio_dqslogic_oct_0}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_4,phy_ddio_dqslogic_readlatency_3,phy_ddio_dqslogic_readlatency_2,phy_ddio_dqslogic_readlatency_1,phy_ddio_dqslogic_readlatency_0}),
	.output_strobe_ena({phy_ddio_dqs_oe_1,phy_ddio_dqs_oe_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_7,phy_ddio_dmdout_6,phy_ddio_dmdout_5,phy_ddio_dmdout_4}),
	.write_data_in({phy_ddio_dqdout_67,phy_ddio_dqdout_66,phy_ddio_dqdout_65,phy_ddio_dqdout_64,phy_ddio_dqdout_63,phy_ddio_dqdout_62,phy_ddio_dqdout_61,phy_ddio_dqdout_60,phy_ddio_dqdout_59,phy_ddio_dqdout_58,phy_ddio_dqdout_57,phy_ddio_dqdout_56,phy_ddio_dqdout_55,phy_ddio_dqdout_54,
phy_ddio_dqdout_53,phy_ddio_dqdout_52,phy_ddio_dqdout_51,phy_ddio_dqdout_50,phy_ddio_dqdout_49,phy_ddio_dqdout_48,phy_ddio_dqdout_47,phy_ddio_dqdout_46,phy_ddio_dqdout_45,phy_ddio_dqdout_44,phy_ddio_dqdout_43,phy_ddio_dqdout_42,phy_ddio_dqdout_41,phy_ddio_dqdout_40,
phy_ddio_dqdout_39,phy_ddio_dqdout_38,phy_ddio_dqdout_37,phy_ddio_dqdout_36}),
	.write_oe_in({phy_ddio_dqoe_33,phy_ddio_dqoe_32,phy_ddio_dqoe_31,phy_ddio_dqoe_30,phy_ddio_dqoe_29,phy_ddio_dqoe_28,phy_ddio_dqoe_27,phy_ddio_dqoe_26,phy_ddio_dqoe_25,phy_ddio_dqoe_24,phy_ddio_dqoe_23,phy_ddio_dqoe_22,phy_ddio_dqoe_21,phy_ddio_dqoe_20,phy_ddio_dqoe_19,phy_ddio_dqoe_18}),
	.write_strobe({phy_ddio_dqs_dout_7,phy_ddio_dqs_dout_6,phy_ddio_dqs_dout_5,phy_ddio_dqs_dout_4}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_1),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_1),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_3,phy_ddio_dqslogic_incrdataen_2}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_3,phy_ddio_dqslogic_incwrptr_2}),
	.oct_ena_in({phy_ddio_dqslogic_oct_3,phy_ddio_dqslogic_oct_2}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_9,phy_ddio_dqslogic_readlatency_8,phy_ddio_dqslogic_readlatency_7,phy_ddio_dqslogic_readlatency_6,phy_ddio_dqslogic_readlatency_5}),
	.output_strobe_ena({phy_ddio_dqs_oe_3,phy_ddio_dqs_oe_2}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_11,phy_ddio_dmdout_10,phy_ddio_dmdout_9,phy_ddio_dmdout_8}),
	.write_data_in({phy_ddio_dqdout_103,phy_ddio_dqdout_102,phy_ddio_dqdout_101,phy_ddio_dqdout_100,phy_ddio_dqdout_99,phy_ddio_dqdout_98,phy_ddio_dqdout_97,phy_ddio_dqdout_96,phy_ddio_dqdout_95,phy_ddio_dqdout_94,phy_ddio_dqdout_93,phy_ddio_dqdout_92,phy_ddio_dqdout_91,phy_ddio_dqdout_90,
phy_ddio_dqdout_89,phy_ddio_dqdout_88,phy_ddio_dqdout_87,phy_ddio_dqdout_86,phy_ddio_dqdout_85,phy_ddio_dqdout_84,phy_ddio_dqdout_83,phy_ddio_dqdout_82,phy_ddio_dqdout_81,phy_ddio_dqdout_80,phy_ddio_dqdout_79,phy_ddio_dqdout_78,phy_ddio_dqdout_77,phy_ddio_dqdout_76,
phy_ddio_dqdout_75,phy_ddio_dqdout_74,phy_ddio_dqdout_73,phy_ddio_dqdout_72}),
	.write_oe_in({phy_ddio_dqoe_51,phy_ddio_dqoe_50,phy_ddio_dqoe_49,phy_ddio_dqoe_48,phy_ddio_dqoe_47,phy_ddio_dqoe_46,phy_ddio_dqoe_45,phy_ddio_dqoe_44,phy_ddio_dqoe_43,phy_ddio_dqoe_42,phy_ddio_dqoe_41,phy_ddio_dqoe_40,phy_ddio_dqoe_39,phy_ddio_dqoe_38,phy_ddio_dqoe_37,phy_ddio_dqoe_36}),
	.write_strobe({phy_ddio_dqs_dout_11,phy_ddio_dqs_dout_10,phy_ddio_dqs_dout_9,phy_ddio_dqs_dout_8}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_2),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_2),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_5,phy_ddio_dqslogic_incrdataen_4}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_5,phy_ddio_dqslogic_incwrptr_4}),
	.oct_ena_in({phy_ddio_dqslogic_oct_5,phy_ddio_dqslogic_oct_4}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_14,phy_ddio_dqslogic_readlatency_13,phy_ddio_dqslogic_readlatency_12,phy_ddio_dqslogic_readlatency_11,phy_ddio_dqslogic_readlatency_10}),
	.output_strobe_ena({phy_ddio_dqs_oe_5,phy_ddio_dqs_oe_4}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_15,phy_ddio_dmdout_14,phy_ddio_dmdout_13,phy_ddio_dmdout_12}),
	.write_data_in({phy_ddio_dqdout_139,phy_ddio_dqdout_138,phy_ddio_dqdout_137,phy_ddio_dqdout_136,phy_ddio_dqdout_135,phy_ddio_dqdout_134,phy_ddio_dqdout_133,phy_ddio_dqdout_132,phy_ddio_dqdout_131,phy_ddio_dqdout_130,phy_ddio_dqdout_129,phy_ddio_dqdout_128,phy_ddio_dqdout_127,
phy_ddio_dqdout_126,phy_ddio_dqdout_125,phy_ddio_dqdout_124,phy_ddio_dqdout_123,phy_ddio_dqdout_122,phy_ddio_dqdout_121,phy_ddio_dqdout_120,phy_ddio_dqdout_119,phy_ddio_dqdout_118,phy_ddio_dqdout_117,phy_ddio_dqdout_116,phy_ddio_dqdout_115,phy_ddio_dqdout_114,
phy_ddio_dqdout_113,phy_ddio_dqdout_112,phy_ddio_dqdout_111,phy_ddio_dqdout_110,phy_ddio_dqdout_109,phy_ddio_dqdout_108}),
	.write_oe_in({phy_ddio_dqoe_69,phy_ddio_dqoe_68,phy_ddio_dqoe_67,phy_ddio_dqoe_66,phy_ddio_dqoe_65,phy_ddio_dqoe_64,phy_ddio_dqoe_63,phy_ddio_dqoe_62,phy_ddio_dqoe_61,phy_ddio_dqoe_60,phy_ddio_dqoe_59,phy_ddio_dqoe_58,phy_ddio_dqoe_57,phy_ddio_dqoe_56,phy_ddio_dqoe_55,phy_ddio_dqoe_54}),
	.write_strobe({phy_ddio_dqs_dout_15,phy_ddio_dqs_dout_14,phy_ddio_dqs_dout_13,phy_ddio_dqs_dout_12}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_3),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_3),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_7,phy_ddio_dqslogic_incrdataen_6}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_7,phy_ddio_dqslogic_incwrptr_6}),
	.oct_ena_in({phy_ddio_dqslogic_oct_7,phy_ddio_dqslogic_oct_6}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_19,phy_ddio_dqslogic_readlatency_18,phy_ddio_dqslogic_readlatency_17,phy_ddio_dqslogic_readlatency_16,phy_ddio_dqslogic_readlatency_15}),
	.output_strobe_ena({phy_ddio_dqs_oe_7,phy_ddio_dqs_oe_6}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_25 (
	pll_dqs_clk,
	pll_hr_clk,
	afi_clk,
	avl_clk,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
input 	pll_hr_clk;
output 	afi_clk;
output 	avl_clk;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;

assign afi_clk = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

assign avl_clk = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(pll_dqs_clk),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_pll (
	pll_mem_clk,
	pll_write_clk)/* synthesis synthesis_greybox=0 */;
output 	pll_mem_clk;
output 	pll_write_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_out[2] ;
wire \clk_out[3] ;

wire [3:0] pll_CLK_OUT_bus;

assign pll_mem_clk = pll_CLK_OUT_bus[0];
assign pll_write_clk = pll_CLK_OUT_bus[1];
assign \clk_out[2]  = pll_CLK_OUT_bus[2];
assign \clk_out[3]  = pll_CLK_OUT_bus[3];

cyclonev_hps_sdram_pll pll(
	.ref_clk(gnd),
	.clk_out(pll_CLK_OUT_bus));

endmodule

module Computer_System_Computer_System_dma_1 (
	f2h_ARREADY_0,
	f2h_RVALID_0,
	outclk_wire_0,
	readaddress_2,
	readaddress_3,
	readaddress_4,
	readaddress_5,
	readaddress_6,
	readaddress_7,
	readaddress_8,
	readaddress_9,
	readaddress_10,
	readaddress_11,
	readaddress_12,
	readaddress_13,
	readaddress_14,
	readaddress_15,
	readaddress_16,
	readaddress_17,
	readaddress_18,
	readaddress_19,
	readaddress_20,
	readaddress_21,
	readaddress_22,
	readaddress_23,
	readaddress_24,
	readaddress_25,
	readaddress_26,
	readaddress_27,
	readaddress_28,
	readaddress_29,
	readaddress_30,
	readaddress_31,
	writeaddress_15,
	q_b_0,
	writeaddress_2,
	writeaddress_3,
	writeaddress_4,
	writeaddress_5,
	writeaddress_6,
	writeaddress_7,
	writeaddress_8,
	writeaddress_9,
	writeaddress_10,
	writeaddress_11,
	writeaddress_12,
	writeaddress_13,
	writeaddress_14,
	writeaddress_1,
	writeaddress_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	mem_used_7,
	saved_grant_0,
	read_select,
	hold_waitrequest,
	write,
	WideOr0,
	wait_latency_counter_1,
	saved_grant_1,
	mem_used_1,
	fifo_empty,
	wren,
	last_write_collision,
	last_write_data_0,
	control_2,
	control_0,
	last_write_data_1,
	last_write_data_2,
	last_write_data_3,
	last_write_data_4,
	last_write_data_5,
	last_write_data_6,
	last_write_data_7,
	write_writedata,
	last_write_data_8,
	write_writedata1,
	last_write_data_9,
	write_writedata2,
	last_write_data_10,
	write_writedata3,
	last_write_data_11,
	write_writedata4,
	last_write_data_12,
	write_writedata5,
	last_write_data_13,
	write_writedata6,
	last_write_data_14,
	write_writedata7,
	last_write_data_15,
	last_write_data_16,
	last_write_data_17,
	last_write_data_18,
	last_write_data_19,
	last_write_data_20,
	last_write_data_21,
	last_write_data_22,
	last_write_data_23,
	last_write_data_24,
	last_write_data_25,
	last_write_data_26,
	last_write_data_27,
	last_write_data_28,
	last_write_data_29,
	last_write_data_30,
	last_write_data_31,
	WideOr1,
	system_reset_n,
	inc_read,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	av_readdatavalid3,
	in_data_reg_2,
	in_data_reg_59,
	mem,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	dma_ctl_readdata_0,
	dma_ctl_readdata_1,
	dma_ctl_readdata_2,
	dma_ctl_readdata_3,
	dma_ctl_readdata_4,
	dma_ctl_readdata_5,
	dma_ctl_readdata_6,
	dma_ctl_readdata_7,
	dma_ctl_readdata_8,
	dma_ctl_readdata_9,
	dma_ctl_readdata_10,
	dma_ctl_readdata_11,
	dma_ctl_readdata_12,
	dma_ctl_readdata_13,
	dma_ctl_readdata_14,
	dma_ctl_readdata_15,
	dma_ctl_readdata_16,
	dma_ctl_readdata_17,
	dma_ctl_readdata_18,
	dma_ctl_readdata_19,
	dma_ctl_readdata_20,
	dma_ctl_readdata_21,
	dma_ctl_readdata_22,
	dma_ctl_readdata_23,
	dma_ctl_readdata_24,
	dma_ctl_readdata_25,
	dma_ctl_readdata_26,
	dma_ctl_readdata_27,
	dma_ctl_readdata_28,
	dma_ctl_readdata_29,
	dma_ctl_readdata_30,
	dma_ctl_readdata_31,
	av_readdatavalid4,
	src0_valid,
	src_data_8,
	src_data_81,
	src_data_16,
	src_data_24,
	src_data_0,
	src_data_01,
	in_data_reg_0,
	in_data_reg_1,
	src_data_9,
	src_data_91,
	src_data_17,
	src_data_25,
	src_data_1,
	src_data_11,
	src_data_10,
	src_data_101,
	src_data_18,
	src_data_26,
	src_data_2,
	src_data_21,
	src_data_111,
	src_data_112,
	src_data_19,
	src_data_27,
	src_data_3,
	src_data_31,
	src_data_12,
	src_data_121,
	src_data_20,
	src_data_28,
	src_data_4,
	src_data_41,
	src_data_13,
	src_data_131,
	src_data_211,
	src_data_29,
	src_data_5,
	src_data_51,
	src_data_14,
	src_data_141,
	src_data_22,
	src_data_30,
	src_data_6,
	src_data_61,
	src_data_15,
	src_data_151,
	src_data_23,
	src_data_311,
	src_data_7,
	src_data_71,
	src_data_82,
	src_data_92,
	src_data_102,
	src_data_113,
	src_data_122,
	src_data_132,
	src_data_142,
	src_data_152)/* synthesis synthesis_greybox=0 */;
input 	f2h_ARREADY_0;
input 	f2h_RVALID_0;
input 	outclk_wire_0;
output 	readaddress_2;
output 	readaddress_3;
output 	readaddress_4;
output 	readaddress_5;
output 	readaddress_6;
output 	readaddress_7;
output 	readaddress_8;
output 	readaddress_9;
output 	readaddress_10;
output 	readaddress_11;
output 	readaddress_12;
output 	readaddress_13;
output 	readaddress_14;
output 	readaddress_15;
output 	readaddress_16;
output 	readaddress_17;
output 	readaddress_18;
output 	readaddress_19;
output 	readaddress_20;
output 	readaddress_21;
output 	readaddress_22;
output 	readaddress_23;
output 	readaddress_24;
output 	readaddress_25;
output 	readaddress_26;
output 	readaddress_27;
output 	readaddress_28;
output 	readaddress_29;
output 	readaddress_30;
output 	readaddress_31;
output 	writeaddress_15;
output 	q_b_0;
output 	writeaddress_2;
output 	writeaddress_3;
output 	writeaddress_4;
output 	writeaddress_5;
output 	writeaddress_6;
output 	writeaddress_7;
output 	writeaddress_8;
output 	writeaddress_9;
output 	writeaddress_10;
output 	writeaddress_11;
output 	writeaddress_12;
output 	writeaddress_13;
output 	writeaddress_14;
output 	writeaddress_1;
output 	writeaddress_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	mem_used_7;
input 	saved_grant_0;
output 	read_select;
input 	hold_waitrequest;
input 	write;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	saved_grant_1;
input 	mem_used_1;
output 	fifo_empty;
input 	wren;
output 	last_write_collision;
output 	last_write_data_0;
output 	control_2;
output 	control_0;
output 	last_write_data_1;
output 	last_write_data_2;
output 	last_write_data_3;
output 	last_write_data_4;
output 	last_write_data_5;
output 	last_write_data_6;
output 	last_write_data_7;
output 	write_writedata;
output 	last_write_data_8;
output 	write_writedata1;
output 	last_write_data_9;
output 	write_writedata2;
output 	last_write_data_10;
output 	write_writedata3;
output 	last_write_data_11;
output 	write_writedata4;
output 	last_write_data_12;
output 	write_writedata5;
output 	last_write_data_13;
output 	write_writedata6;
output 	last_write_data_14;
output 	write_writedata7;
output 	last_write_data_15;
output 	last_write_data_16;
output 	last_write_data_17;
output 	last_write_data_18;
output 	last_write_data_19;
output 	last_write_data_20;
output 	last_write_data_21;
output 	last_write_data_22;
output 	last_write_data_23;
output 	last_write_data_24;
output 	last_write_data_25;
output 	last_write_data_26;
output 	last_write_data_27;
output 	last_write_data_28;
output 	last_write_data_29;
output 	last_write_data_30;
output 	last_write_data_31;
input 	WideOr1;
input 	system_reset_n;
output 	inc_read;
input 	av_readdatavalid;
input 	av_readdatavalid1;
input 	av_readdatavalid2;
input 	av_readdatavalid3;
input 	in_data_reg_2;
input 	in_data_reg_59;
input 	mem;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_4;
input 	int_nxt_addr_reg_dly_3;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
output 	dma_ctl_readdata_0;
output 	dma_ctl_readdata_1;
output 	dma_ctl_readdata_2;
output 	dma_ctl_readdata_3;
output 	dma_ctl_readdata_4;
output 	dma_ctl_readdata_5;
output 	dma_ctl_readdata_6;
output 	dma_ctl_readdata_7;
output 	dma_ctl_readdata_8;
output 	dma_ctl_readdata_9;
output 	dma_ctl_readdata_10;
output 	dma_ctl_readdata_11;
output 	dma_ctl_readdata_12;
output 	dma_ctl_readdata_13;
output 	dma_ctl_readdata_14;
output 	dma_ctl_readdata_15;
output 	dma_ctl_readdata_16;
output 	dma_ctl_readdata_17;
output 	dma_ctl_readdata_18;
output 	dma_ctl_readdata_19;
output 	dma_ctl_readdata_20;
output 	dma_ctl_readdata_21;
output 	dma_ctl_readdata_22;
output 	dma_ctl_readdata_23;
output 	dma_ctl_readdata_24;
output 	dma_ctl_readdata_25;
output 	dma_ctl_readdata_26;
output 	dma_ctl_readdata_27;
output 	dma_ctl_readdata_28;
output 	dma_ctl_readdata_29;
output 	dma_ctl_readdata_30;
output 	dma_ctl_readdata_31;
input 	av_readdatavalid4;
input 	src0_valid;
input 	src_data_8;
input 	src_data_81;
input 	src_data_16;
input 	src_data_24;
input 	src_data_0;
input 	src_data_01;
input 	in_data_reg_0;
input 	in_data_reg_1;
input 	src_data_9;
input 	src_data_91;
input 	src_data_17;
input 	src_data_25;
input 	src_data_1;
input 	src_data_11;
input 	src_data_10;
input 	src_data_101;
input 	src_data_18;
input 	src_data_26;
input 	src_data_2;
input 	src_data_21;
input 	src_data_111;
input 	src_data_112;
input 	src_data_19;
input 	src_data_27;
input 	src_data_3;
input 	src_data_31;
input 	src_data_12;
input 	src_data_121;
input 	src_data_20;
input 	src_data_28;
input 	src_data_4;
input 	src_data_41;
input 	src_data_13;
input 	src_data_131;
input 	src_data_211;
input 	src_data_29;
input 	src_data_5;
input 	src_data_51;
input 	src_data_14;
input 	src_data_141;
input 	src_data_22;
input 	src_data_30;
input 	src_data_6;
input 	src_data_61;
input 	src_data_15;
input 	src_data_151;
input 	src_data_23;
input 	src_data_311;
input 	src_data_7;
input 	src_data_71;
input 	src_data_82;
input 	src_data_92;
input 	src_data_102;
input 	src_data_113;
input 	src_data_122;
input 	src_data_132;
input 	src_data_142;
input 	src_data_152;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add2~1_sumout ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add2~7 ;
wire \Add2~9_sumout ;
wire \Add2~10 ;
wire \Add2~11 ;
wire \Add2~13_sumout ;
wire \Add2~14 ;
wire \Add2~15 ;
wire \Add2~17_sumout ;
wire \Add2~18 ;
wire \Add2~19 ;
wire \Add2~21_sumout ;
wire \Add2~22 ;
wire \Add2~23 ;
wire \Add2~25_sumout ;
wire \Add2~26 ;
wire \Add2~27 ;
wire \Add2~29_sumout ;
wire \Add2~30 ;
wire \Add2~31 ;
wire \Add2~33_sumout ;
wire \Add2~34 ;
wire \Add2~35 ;
wire \Add2~37_sumout ;
wire \Add2~38 ;
wire \Add2~39 ;
wire \Add2~41_sumout ;
wire \Add2~42 ;
wire \Add2~43 ;
wire \Add2~45_sumout ;
wire \Add2~46 ;
wire \Add2~47 ;
wire \Add2~49_sumout ;
wire \Add2~50 ;
wire \Add2~51 ;
wire \Add2~53_sumout ;
wire \Add2~54 ;
wire \Add2~55 ;
wire \Add2~57_sumout ;
wire \Add2~58 ;
wire \Add2~59 ;
wire \Add2~61_sumout ;
wire \Add2~62 ;
wire \Add2~63 ;
wire \Add2~65_sumout ;
wire \Add2~66 ;
wire \Add2~67 ;
wire \Add2~69_sumout ;
wire \Add2~70 ;
wire \Add2~71 ;
wire \Add2~73_sumout ;
wire \Add2~74 ;
wire \Add2~75 ;
wire \Add2~77_sumout ;
wire \Add2~78 ;
wire \Add2~79 ;
wire \Add2~81_sumout ;
wire \Add2~82 ;
wire \Add2~83 ;
wire \Add2~85_sumout ;
wire \Add2~86 ;
wire \Add2~87 ;
wire \Add2~89_sumout ;
wire \Add2~90 ;
wire \Add2~91 ;
wire \Add2~93_sumout ;
wire \Add2~94 ;
wire \Add2~95 ;
wire \Add2~97_sumout ;
wire \Add2~98 ;
wire \Add2~99 ;
wire \Add2~101_sumout ;
wire \Add2~102 ;
wire \Add2~103 ;
wire \Add2~105_sumout ;
wire \Add2~106 ;
wire \Add2~107 ;
wire \Add2~109_sumout ;
wire \Add2~110 ;
wire \Add2~111 ;
wire \Add2~113_sumout ;
wire \Add2~114 ;
wire \Add2~115 ;
wire \Add2~117_sumout ;
wire \Add2~118 ;
wire \Add2~119 ;
wire \Add2~121_sumout ;
wire \Add2~122 ;
wire \Add2~123 ;
wire \Add2~125_sumout ;
wire \Add2~126 ;
wire \Add2~127 ;
wire \length[31]~q ;
wire \length[22]~q ;
wire \length[23]~q ;
wire \length[24]~q ;
wire \length[25]~q ;
wire \length[26]~q ;
wire \length[12]~q ;
wire \length[13]~q ;
wire \length[14]~q ;
wire \length[15]~q ;
wire \length[16]~q ;
wire \length[1]~q ;
wire \length[2]~q ;
wire \length[3]~q ;
wire \length[4]~q ;
wire \length[5]~q ;
wire \length[6]~q ;
wire \length[27]~q ;
wire \length[28]~q ;
wire \length[29]~q ;
wire \length[11]~q ;
wire \length[20]~q ;
wire \length[21]~q ;
wire \length[30]~q ;
wire \length[17]~q ;
wire \length[18]~q ;
wire \length[19]~q ;
wire \length[0]~q ;
wire \length[7]~q ;
wire \length[8]~q ;
wire \length[9]~q ;
wire \length[10]~q ;
wire \p1_writelength_eq_0~0_combout ;
wire \p1_writelength_eq_0~1_combout ;
wire \p1_writelength_eq_0~2_combout ;
wire \p1_done_write~0_combout ;
wire \length_eq_0~q ;
wire \p1_length_eq_0~0_combout ;
wire \p1_length_eq_0~1_combout ;
wire \p1_length_eq_0~2_combout ;
wire \p1_length_eq_0~3_combout ;
wire \p1_length_eq_0~4_combout ;
wire \p1_length_eq_0~5_combout ;
wire \p1_length_eq_0~6_combout ;
wire \p1_length_eq_0~7_combout ;
wire \p1_done_read~0_combout ;
wire \the_Computer_System_dma_1_fifo_module|p1_fifo_full~3_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[0]~3_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[1]~6_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[2]~9_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[3]~12_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[4]~15_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[5]~18_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[6]~21_combout ;
wire \the_Computer_System_dma_1_read_data_mux|fifo_wr_data[7]~24_combout ;
wire \length_eq_0~0_combout ;
wire \length[29]~0_combout ;
wire \p1_readaddress~1_combout ;
wire \Equal3~2_combout ;
wire \p1_control~0_combout ;
wire \control[12]~q ;
wire \set_software_reset_bit~0_combout ;
wire \d1_softwarereset~0_combout ;
wire \d1_softwarereset~q ;
wire \software_reset_request~0_combout ;
wire \software_reset_request~q ;
wire \reset_n~0_combout ;
wire \reset_n~q ;
wire \control[8]~q ;
wire \Add0~125_sumout ;
wire \Equal3~0_combout ;
wire \p1_readaddress~0_combout ;
wire \readaddress[27]~0_combout ;
wire \readaddress[0]~q ;
wire \Add0~126 ;
wire \Add0~121_sumout ;
wire \readaddress[1]~q ;
wire \Add0~122 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \Add0~110 ;
wire \Add0~113_sumout ;
wire \Add0~114 ;
wire \Add0~117_sumout ;
wire \control[9]~q ;
wire \Add1~62 ;
wire \Add1~58 ;
wire \Add1~6 ;
wire \Add1~10 ;
wire \Add1~14 ;
wire \Add1~18 ;
wire \Add1~22 ;
wire \Add1~26 ;
wire \Add1~30 ;
wire \Add1~34 ;
wire \Add1~38 ;
wire \Add1~42 ;
wire \Add1~46 ;
wire \Add1~50 ;
wire \Add1~54 ;
wire \Add1~1_sumout ;
wire \Equal3~1_combout ;
wire \p1_writeaddress~0_combout ;
wire \writeaddress[8]~0_combout ;
wire \Add1~5_sumout ;
wire \Add1~9_sumout ;
wire \Add1~13_sumout ;
wire \Add1~17_sumout ;
wire \Add1~21_sumout ;
wire \Add1~25_sumout ;
wire \Add1~29_sumout ;
wire \Add1~33_sumout ;
wire \Add1~37_sumout ;
wire \Add1~41_sumout ;
wire \Add1~45_sumout ;
wire \Add1~49_sumout ;
wire \Add1~53_sumout ;
wire \Add1~57_sumout ;
wire \Add1~61_sumout ;
wire \control[2]~0_combout ;
wire \Add3~109_sumout ;
wire \Equal3~3_combout ;
wire \p1_length~0_combout ;
wire \writelength[30]~q ;
wire \Add3~110 ;
wire \Add3~111 ;
wire \Add3~113_sumout ;
wire \writelength[1]~q ;
wire \Add3~114 ;
wire \Add3~115 ;
wire \Add3~117_sumout ;
wire \writelength[2]~q ;
wire \Add3~118 ;
wire \Add3~119 ;
wire \Add3~121_sumout ;
wire \writelength[3]~q ;
wire \Add3~122 ;
wire \Add3~123 ;
wire \Add3~125_sumout ;
wire \writelength[4]~q ;
wire \Add3~126 ;
wire \Add3~127 ;
wire \Add3~53_sumout ;
wire \writelength[5]~q ;
wire \Add3~54 ;
wire \Add3~55 ;
wire \Add3~57_sumout ;
wire \writelength[6]~q ;
wire \Add3~58 ;
wire \Add3~59 ;
wire \Add3~61_sumout ;
wire \writelength[7]~q ;
wire \Add3~62 ;
wire \Add3~63 ;
wire \Add3~65_sumout ;
wire \writelength[8]~q ;
wire \Add3~66 ;
wire \Add3~67 ;
wire \Add3~33_sumout ;
wire \writelength[9]~q ;
wire \Add3~34 ;
wire \Add3~35 ;
wire \Add3~89_sumout ;
wire \writelength[10]~q ;
wire \Add3~90 ;
wire \Add3~91 ;
wire \Add3~93_sumout ;
wire \writelength[11]~q ;
wire \Add3~94 ;
wire \Add3~95 ;
wire \Add3~97_sumout ;
wire \writelength[12]~q ;
wire \Add3~98 ;
wire \Add3~99 ;
wire \Add3~101_sumout ;
wire \writelength[13]~q ;
wire \Add3~102 ;
wire \Add3~103 ;
wire \Add3~37_sumout ;
wire \writelength[14]~q ;
wire \Add3~38 ;
wire \Add3~39 ;
wire \Add3~105_sumout ;
wire \writelength[15]~q ;
wire \Add3~106 ;
wire \Add3~107 ;
wire \Add3~41_sumout ;
wire \writelength[16]~q ;
wire \Add3~42 ;
wire \Add3~43 ;
wire \Add3~45_sumout ;
wire \writelength[17]~q ;
wire \Add3~46 ;
wire \Add3~47 ;
wire \Add3~49_sumout ;
wire \writelength[18]~q ;
wire \Add3~50 ;
wire \Add3~51 ;
wire \Add3~13_sumout ;
wire \writelength[19]~q ;
wire \Add3~14 ;
wire \Add3~15 ;
wire \Add3~69_sumout ;
wire \writelength[20]~q ;
wire \Add3~70 ;
wire \Add3~71 ;
wire \Add3~73_sumout ;
wire \writelength[21]~q ;
wire \Add3~74 ;
wire \Add3~75 ;
wire \Add3~77_sumout ;
wire \writelength[22]~q ;
wire \Add3~78 ;
wire \Add3~79 ;
wire \Add3~81_sumout ;
wire \writelength[23]~q ;
wire \Add3~82 ;
wire \Add3~83 ;
wire \Add3~17_sumout ;
wire \writelength[24]~q ;
wire \Add3~18 ;
wire \Add3~19 ;
wire \Add3~85_sumout ;
wire \writelength[25]~q ;
wire \Add3~86 ;
wire \Add3~87 ;
wire \Add3~21_sumout ;
wire \writelength[26]~q ;
wire \Add3~22 ;
wire \Add3~23 ;
wire \Add3~25_sumout ;
wire \writelength[27]~q ;
wire \Add3~26 ;
wire \Add3~27 ;
wire \Add3~29_sumout ;
wire \writelength[28]~q ;
wire \Add3~30 ;
wire \Add3~31 ;
wire \Add3~1_sumout ;
wire \writelength[29]~q ;
wire \Add3~2 ;
wire \Add3~3 ;
wire \Add3~5_sumout ;
wire \writelength[31]~q ;
wire \Add3~6 ;
wire \Add3~7 ;
wire \Add3~9_sumout ;
wire \p1_writelength_eq_0~6_combout ;
wire \p1_writelength_eq_0~7_combout ;
wire \p1_writelength_eq_0~8_combout ;
wire \p1_writelength_eq_0~3_combout ;
wire \p1_writelength_eq_0~4_combout ;
wire \p1_writelength_eq_0~5_combout ;
wire \writelength_eq_0~0_combout ;
wire \writelength_eq_0~q ;
wire \writelength[13]~0_combout ;
wire \writelength[13]~1_combout ;
wire \writelength[0]~q ;
wire \p1_dma_ctl_readdata[0]~0_combout ;
wire \Equal3~4_combout ;
wire \control[3]~q ;
wire \control[7]~1_combout ;
wire \control[7]~q ;
wire \p1_done_write~1_combout ;
wire \done_write~q ;
wire \done_transaction~combout ;
wire \d1_done_transaction~q ;
wire \flush_fifo~combout ;
wire \p1_dma_ctl_readdata~1_combout ;
wire \done~0_combout ;
wire \done~q ;
wire \p1_dma_ctl_readdata[0]~2_combout ;
wire \p1_dma_ctl_readdata[0]~combout ;
wire \p1_dma_ctl_readdata[1]~3_combout ;
wire \control[1]~q ;
wire \p1_dma_ctl_readdata[1]~4_combout ;
wire \p1_dma_ctl_readdata[1]~combout ;
wire \p1_dma_ctl_readdata[2]~43_combout ;
wire \p1_dma_ctl_readdata[3]~39_combout ;
wire \p1_dma_ctl_readdata[4]~5_combout ;
wire \control[4]~q ;
wire \len~0_combout ;
wire \len~q ;
wire \p1_dma_ctl_readdata[4]~6_combout ;
wire \p1_dma_ctl_readdata[4]~combout ;
wire \control[5]~q ;
wire \p1_dma_ctl_readdata[5]~35_combout ;
wire \control[6]~q ;
wire \p1_dma_ctl_readdata[6]~31_combout ;
wire \p1_dma_ctl_readdata[7]~27_combout ;
wire \p1_dma_ctl_readdata[8]~23_combout ;
wire \p1_dma_ctl_readdata[9]~19_combout ;
wire \control[10]~q ;
wire \p1_dma_ctl_readdata[10]~15_combout ;
wire \control[11]~q ;
wire \p1_dma_ctl_readdata[11]~11_combout ;
wire \p1_dma_ctl_readdata[12]~7_combout ;
wire \p1_dma_ctl_readdata[13]~combout ;
wire \p1_dma_ctl_readdata[14]~combout ;
wire \p1_dma_ctl_readdata[15]~combout ;
wire \Add1~2 ;
wire \Add1~65_sumout ;
wire \writeaddress[16]~q ;
wire \p1_dma_ctl_readdata[16]~combout ;
wire \Add1~66 ;
wire \Add1~69_sumout ;
wire \writeaddress[17]~q ;
wire \p1_dma_ctl_readdata[17]~combout ;
wire \Add1~70 ;
wire \Add1~73_sumout ;
wire \writeaddress[18]~q ;
wire \p1_dma_ctl_readdata[18]~combout ;
wire \Add1~74 ;
wire \Add1~77_sumout ;
wire \writeaddress[19]~q ;
wire \p1_dma_ctl_readdata[19]~combout ;
wire \Add1~78 ;
wire \Add1~81_sumout ;
wire \writeaddress[20]~q ;
wire \p1_dma_ctl_readdata[20]~combout ;
wire \Add1~82 ;
wire \Add1~85_sumout ;
wire \writeaddress[21]~q ;
wire \p1_dma_ctl_readdata[21]~combout ;
wire \Add1~86 ;
wire \Add1~89_sumout ;
wire \writeaddress[22]~q ;
wire \p1_dma_ctl_readdata[22]~combout ;
wire \Add1~90 ;
wire \Add1~93_sumout ;
wire \writeaddress[23]~q ;
wire \p1_dma_ctl_readdata[23]~combout ;
wire \Add1~94 ;
wire \Add1~97_sumout ;
wire \writeaddress[24]~q ;
wire \p1_dma_ctl_readdata[24]~combout ;
wire \Add1~98 ;
wire \Add1~101_sumout ;
wire \writeaddress[25]~q ;
wire \p1_dma_ctl_readdata[25]~combout ;
wire \Add1~102 ;
wire \Add1~105_sumout ;
wire \writeaddress[26]~q ;
wire \p1_dma_ctl_readdata[26]~combout ;
wire \Add1~106 ;
wire \Add1~109_sumout ;
wire \writeaddress[27]~q ;
wire \p1_dma_ctl_readdata[27]~combout ;
wire \p1_dma_ctl_readdata[28]~combout ;
wire \p1_dma_ctl_readdata[29]~combout ;
wire \p1_dma_ctl_readdata[30]~combout ;
wire \p1_dma_ctl_readdata[31]~combout ;


Computer_System_Computer_System_dma_1_mem_read the_Computer_System_dma_1_mem_read(
	.f2h_ARREADY_0(f2h_ARREADY_0),
	.clk(outclk_wire_0),
	.mem_used_7(mem_used_7),
	.saved_grant_0(saved_grant_0),
	.read_select1(read_select),
	.hold_waitrequest(hold_waitrequest),
	.write(write),
	.WideOr1(WideOr1),
	.inc_read1(inc_read),
	.control_3(\control[3]~q ),
	.control_7(\control[7]~q ),
	.p1_done_write(\p1_done_write~0_combout ),
	.p1_done_read(\p1_done_read~0_combout ),
	.p1_fifo_full(\the_Computer_System_dma_1_fifo_module|p1_fifo_full~3_combout ),
	.reset_n(\reset_n~q ));

Computer_System_Computer_System_dma_1_fifo_module the_Computer_System_dma_1_fifo_module(
	.outclk_wire_0(outclk_wire_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.fifo_empty1(fifo_empty),
	.wren(wren),
	.last_write_collision1(last_write_collision),
	.last_write_data_0(last_write_data_0),
	.last_write_data_1(last_write_data_1),
	.last_write_data_2(last_write_data_2),
	.last_write_data_3(last_write_data_3),
	.last_write_data_4(last_write_data_4),
	.last_write_data_5(last_write_data_5),
	.last_write_data_6(last_write_data_6),
	.last_write_data_7(last_write_data_7),
	.last_write_data_8(last_write_data_8),
	.last_write_data_9(last_write_data_9),
	.last_write_data_10(last_write_data_10),
	.last_write_data_11(last_write_data_11),
	.last_write_data_12(last_write_data_12),
	.last_write_data_13(last_write_data_13),
	.last_write_data_14(last_write_data_14),
	.last_write_data_15(last_write_data_15),
	.last_write_data_16(last_write_data_16),
	.last_write_data_17(last_write_data_17),
	.last_write_data_18(last_write_data_18),
	.last_write_data_19(last_write_data_19),
	.last_write_data_20(last_write_data_20),
	.last_write_data_21(last_write_data_21),
	.last_write_data_22(last_write_data_22),
	.last_write_data_23(last_write_data_23),
	.last_write_data_24(last_write_data_24),
	.last_write_data_25(last_write_data_25),
	.last_write_data_26(last_write_data_26),
	.last_write_data_27(last_write_data_27),
	.last_write_data_28(last_write_data_28),
	.last_write_data_29(last_write_data_29),
	.last_write_data_30(last_write_data_30),
	.last_write_data_31(last_write_data_31),
	.inc_read(inc_read),
	.flush_fifo(\flush_fifo~combout ),
	.av_readdatavalid(av_readdatavalid),
	.av_readdatavalid1(av_readdatavalid1),
	.av_readdatavalid2(av_readdatavalid2),
	.av_readdatavalid3(av_readdatavalid3),
	.p1_fifo_full(\the_Computer_System_dma_1_fifo_module|p1_fifo_full~3_combout ),
	.reset_n(\reset_n~q ),
	.av_readdatavalid4(av_readdatavalid4),
	.src0_valid(src0_valid),
	.src_data_16(src_data_16),
	.src_data_24(src_data_24),
	.fifo_wr_data_0(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[0]~3_combout ),
	.src_data_17(src_data_17),
	.src_data_25(src_data_25),
	.fifo_wr_data_1(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[1]~6_combout ),
	.src_data_18(src_data_18),
	.src_data_26(src_data_26),
	.fifo_wr_data_2(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[2]~9_combout ),
	.src_data_19(src_data_19),
	.src_data_27(src_data_27),
	.fifo_wr_data_3(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[3]~12_combout ),
	.src_data_20(src_data_20),
	.src_data_28(src_data_28),
	.fifo_wr_data_4(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[4]~15_combout ),
	.src_data_21(src_data_211),
	.src_data_29(src_data_29),
	.fifo_wr_data_5(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[5]~18_combout ),
	.src_data_22(src_data_22),
	.src_data_30(src_data_30),
	.fifo_wr_data_6(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[6]~21_combout ),
	.src_data_23(src_data_23),
	.src_data_31(src_data_311),
	.fifo_wr_data_7(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[7]~24_combout ),
	.src_data_8(src_data_82),
	.src_data_9(src_data_92),
	.src_data_10(src_data_102),
	.src_data_11(src_data_113),
	.src_data_12(src_data_122),
	.src_data_13(src_data_132),
	.src_data_14(src_data_142),
	.src_data_15(src_data_152));

Computer_System_Computer_System_dma_1_read_data_mux the_Computer_System_dma_1_read_data_mux(
	.f2h_RVALID_0(f2h_RVALID_0),
	.clk(outclk_wire_0),
	.readaddress_0(\readaddress[0]~q ),
	.readaddress_1(\readaddress[1]~q ),
	.WideOr0(WideOr0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.control_2(control_2),
	.control_0(control_0),
	.av_readdatavalid(av_readdatavalid),
	.av_readdatavalid1(av_readdatavalid1),
	.av_readdatavalid2(av_readdatavalid2),
	.reset_n(\reset_n~q ),
	.in_data_reg_59(in_data_reg_59),
	.mem(mem),
	.in_data_reg_3(in_data_reg_3),
	.src0_valid(src0_valid),
	.src_data_8(src_data_8),
	.src_data_81(src_data_81),
	.src_data_16(src_data_16),
	.src_data_24(src_data_24),
	.src_data_0(src_data_0),
	.src_data_01(src_data_01),
	.fifo_wr_data_0(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[0]~3_combout ),
	.Equal3(\Equal3~2_combout ),
	.src_data_9(src_data_9),
	.src_data_91(src_data_91),
	.src_data_17(src_data_17),
	.src_data_25(src_data_25),
	.src_data_1(src_data_1),
	.src_data_11(src_data_11),
	.fifo_wr_data_1(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[1]~6_combout ),
	.src_data_10(src_data_10),
	.src_data_101(src_data_101),
	.src_data_18(src_data_18),
	.src_data_26(src_data_26),
	.src_data_2(src_data_2),
	.src_data_21(src_data_21),
	.fifo_wr_data_2(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[2]~9_combout ),
	.src_data_111(src_data_111),
	.src_data_112(src_data_112),
	.src_data_19(src_data_19),
	.src_data_27(src_data_27),
	.src_data_3(src_data_3),
	.src_data_31(src_data_31),
	.fifo_wr_data_3(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[3]~12_combout ),
	.src_data_12(src_data_12),
	.src_data_121(src_data_121),
	.src_data_20(src_data_20),
	.src_data_28(src_data_28),
	.src_data_4(src_data_4),
	.src_data_41(src_data_41),
	.fifo_wr_data_4(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[4]~15_combout ),
	.src_data_13(src_data_13),
	.src_data_131(src_data_131),
	.src_data_211(src_data_211),
	.src_data_29(src_data_29),
	.src_data_5(src_data_5),
	.src_data_51(src_data_51),
	.fifo_wr_data_5(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[5]~18_combout ),
	.src_data_14(src_data_14),
	.src_data_141(src_data_141),
	.src_data_22(src_data_22),
	.src_data_30(src_data_30),
	.src_data_6(src_data_6),
	.src_data_61(src_data_61),
	.fifo_wr_data_6(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[6]~21_combout ),
	.src_data_15(src_data_15),
	.src_data_151(src_data_151),
	.src_data_23(src_data_23),
	.src_data_311(src_data_311),
	.src_data_7(src_data_7),
	.src_data_71(src_data_71),
	.fifo_wr_data_7(\the_Computer_System_dma_1_read_data_mux|fifo_wr_data[7]~24_combout ),
	.p1_length(\p1_length~0_combout ),
	.control_8(\control[8]~q ));

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~94 ),
	.sharein(\Add2~95 ),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h000000000000FF00;
defparam \Add2~1 .shared_arith = "on";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~90 ),
	.sharein(\Add2~91 ),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout(\Add2~7 ));
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~5 .shared_arith = "on";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(\Add2~7 ),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout(\Add2~11 ));
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~9 .shared_arith = "on";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(\Add2~11 ),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout(\Add2~15 ));
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~13 .shared_arith = "on";

cyclonev_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(\Add2~15 ),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout(\Add2~19 ));
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~17 .shared_arith = "on";

cyclonev_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(\Add2~19 ),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout(\Add2~23 ));
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~21 .shared_arith = "on";

cyclonev_lcell_comb \Add2~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~82 ),
	.sharein(\Add2~83 ),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(\Add2~26 ),
	.shareout(\Add2~27 ));
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~25 .shared_arith = "on";

cyclonev_lcell_comb \Add2~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~26 ),
	.sharein(\Add2~27 ),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout(\Add2~31 ));
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~29 .shared_arith = "on";

cyclonev_lcell_comb \Add2~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(\Add2~31 ),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout(\Add2~35 ));
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~33 .shared_arith = "on";

cyclonev_lcell_comb \Add2~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(\Add2~35 ),
	.combout(),
	.sumout(\Add2~37_sumout ),
	.cout(\Add2~38 ),
	.shareout(\Add2~39 ));
defparam \Add2~37 .extended_lut = "off";
defparam \Add2~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~37 .shared_arith = "on";

cyclonev_lcell_comb \Add2~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~38 ),
	.sharein(\Add2~39 ),
	.combout(),
	.sumout(\Add2~41_sumout ),
	.cout(\Add2~42 ),
	.shareout(\Add2~43 ));
defparam \Add2~41 .extended_lut = "off";
defparam \Add2~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~41 .shared_arith = "on";

cyclonev_lcell_comb \Add2~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~110 ),
	.sharein(\Add2~111 ),
	.combout(),
	.sumout(\Add2~45_sumout ),
	.cout(\Add2~46 ),
	.shareout(\Add2~47 ));
defparam \Add2~45 .extended_lut = "off";
defparam \Add2~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~45 .shared_arith = "on";

cyclonev_lcell_comb \Add2~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_2),
	.datad(!\length[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~46 ),
	.sharein(\Add2~47 ),
	.combout(),
	.sumout(\Add2~49_sumout ),
	.cout(\Add2~50 ),
	.shareout(\Add2~51 ));
defparam \Add2~49 .extended_lut = "off";
defparam \Add2~49 .lut_mask = 64'h0000000F00000FF0;
defparam \Add2~49 .shared_arith = "on";

cyclonev_lcell_comb \Add2~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~50 ),
	.sharein(\Add2~51 ),
	.combout(),
	.sumout(\Add2~53_sumout ),
	.cout(\Add2~54 ),
	.shareout(\Add2~55 ));
defparam \Add2~53 .extended_lut = "off";
defparam \Add2~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~53 .shared_arith = "on";

cyclonev_lcell_comb \Add2~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~54 ),
	.sharein(\Add2~55 ),
	.combout(),
	.sumout(\Add2~57_sumout ),
	.cout(\Add2~58 ),
	.shareout(\Add2~59 ));
defparam \Add2~57 .extended_lut = "off";
defparam \Add2~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~57 .shared_arith = "on";

cyclonev_lcell_comb \Add2~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~58 ),
	.sharein(\Add2~59 ),
	.combout(),
	.sumout(\Add2~61_sumout ),
	.cout(\Add2~62 ),
	.shareout(\Add2~63 ));
defparam \Add2~61 .extended_lut = "off";
defparam \Add2~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~61 .shared_arith = "on";

cyclonev_lcell_comb \Add2~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~62 ),
	.sharein(\Add2~63 ),
	.combout(),
	.sumout(\Add2~65_sumout ),
	.cout(\Add2~66 ),
	.shareout(\Add2~67 ));
defparam \Add2~65 .extended_lut = "off";
defparam \Add2~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~65 .shared_arith = "on";

cyclonev_lcell_comb \Add2~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(\Add2~23 ),
	.combout(),
	.sumout(\Add2~69_sumout ),
	.cout(\Add2~70 ),
	.shareout(\Add2~71 ));
defparam \Add2~69 .extended_lut = "off";
defparam \Add2~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~69 .shared_arith = "on";

cyclonev_lcell_comb \Add2~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~70 ),
	.sharein(\Add2~71 ),
	.combout(),
	.sumout(\Add2~73_sumout ),
	.cout(\Add2~74 ),
	.shareout(\Add2~75 ));
defparam \Add2~73 .extended_lut = "off";
defparam \Add2~73 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~73 .shared_arith = "on";

cyclonev_lcell_comb \Add2~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~74 ),
	.sharein(\Add2~75 ),
	.combout(),
	.sumout(\Add2~77_sumout ),
	.cout(\Add2~78 ),
	.shareout(\Add2~79 ));
defparam \Add2~77 .extended_lut = "off";
defparam \Add2~77 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~77 .shared_arith = "on";

cyclonev_lcell_comb \Add2~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~126 ),
	.sharein(\Add2~127 ),
	.combout(),
	.sumout(\Add2~81_sumout ),
	.cout(\Add2~82 ),
	.shareout(\Add2~83 ));
defparam \Add2~81 .extended_lut = "off";
defparam \Add2~81 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~81 .shared_arith = "on";

cyclonev_lcell_comb \Add2~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~106 ),
	.sharein(\Add2~107 ),
	.combout(),
	.sumout(\Add2~85_sumout ),
	.cout(\Add2~86 ),
	.shareout(\Add2~87 ));
defparam \Add2~85 .extended_lut = "off";
defparam \Add2~85 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~85 .shared_arith = "on";

cyclonev_lcell_comb \Add2~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~86 ),
	.sharein(\Add2~87 ),
	.combout(),
	.sumout(\Add2~89_sumout ),
	.cout(\Add2~90 ),
	.shareout(\Add2~91 ));
defparam \Add2~89 .extended_lut = "off";
defparam \Add2~89 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~89 .shared_arith = "on";

cyclonev_lcell_comb \Add2~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~78 ),
	.sharein(\Add2~79 ),
	.combout(),
	.sumout(\Add2~93_sumout ),
	.cout(\Add2~94 ),
	.shareout(\Add2~95 ));
defparam \Add2~93 .extended_lut = "off";
defparam \Add2~93 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~93 .shared_arith = "on";

cyclonev_lcell_comb \Add2~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~42 ),
	.sharein(\Add2~43 ),
	.combout(),
	.sumout(\Add2~97_sumout ),
	.cout(\Add2~98 ),
	.shareout(\Add2~99 ));
defparam \Add2~97 .extended_lut = "off";
defparam \Add2~97 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~97 .shared_arith = "on";

cyclonev_lcell_comb \Add2~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~98 ),
	.sharein(\Add2~99 ),
	.combout(),
	.sumout(\Add2~101_sumout ),
	.cout(\Add2~102 ),
	.shareout(\Add2~103 ));
defparam \Add2~101 .extended_lut = "off";
defparam \Add2~101 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~101 .shared_arith = "on";

cyclonev_lcell_comb \Add2~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~102 ),
	.sharein(\Add2~103 ),
	.combout(),
	.sumout(\Add2~105_sumout ),
	.cout(\Add2~106 ),
	.shareout(\Add2~107 ));
defparam \Add2~105 .extended_lut = "off";
defparam \Add2~105 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~105 .shared_arith = "on";

cyclonev_lcell_comb \Add2~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_0),
	.datad(!\length[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~109_sumout ),
	.cout(\Add2~110 ),
	.shareout(\Add2~111 ));
defparam \Add2~109 .extended_lut = "off";
defparam \Add2~109 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~109 .shared_arith = "on";

cyclonev_lcell_comb \Add2~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~66 ),
	.sharein(\Add2~67 ),
	.combout(),
	.sumout(\Add2~113_sumout ),
	.cout(\Add2~114 ),
	.shareout(\Add2~115 ));
defparam \Add2~113 .extended_lut = "off";
defparam \Add2~113 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~113 .shared_arith = "on";

cyclonev_lcell_comb \Add2~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~114 ),
	.sharein(\Add2~115 ),
	.combout(),
	.sumout(\Add2~117_sumout ),
	.cout(\Add2~118 ),
	.shareout(\Add2~119 ));
defparam \Add2~117 .extended_lut = "off";
defparam \Add2~117 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~117 .shared_arith = "on";

cyclonev_lcell_comb \Add2~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~118 ),
	.sharein(\Add2~119 ),
	.combout(),
	.sumout(\Add2~121_sumout ),
	.cout(\Add2~122 ),
	.shareout(\Add2~123 ));
defparam \Add2~121 .extended_lut = "off";
defparam \Add2~121 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~121 .shared_arith = "on";

cyclonev_lcell_comb \Add2~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~122 ),
	.sharein(\Add2~123 ),
	.combout(),
	.sumout(\Add2~125_sumout ),
	.cout(\Add2~126 ),
	.shareout(\Add2~127 ));
defparam \Add2~125 .extended_lut = "off";
defparam \Add2~125 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~125 .shared_arith = "on";

dffeas \length[31] (
	.clk(outclk_wire_0),
	.d(in_data_reg_31),
	.asdata(\Add2~1_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[31]~q ),
	.prn(vcc));
defparam \length[31] .is_wysiwyg = "true";
defparam \length[31] .power_up = "low";

dffeas \length[22] (
	.clk(outclk_wire_0),
	.d(in_data_reg_22),
	.asdata(\Add2~5_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[22]~q ),
	.prn(vcc));
defparam \length[22] .is_wysiwyg = "true";
defparam \length[22] .power_up = "low";

dffeas \length[23] (
	.clk(outclk_wire_0),
	.d(in_data_reg_23),
	.asdata(\Add2~9_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[23]~q ),
	.prn(vcc));
defparam \length[23] .is_wysiwyg = "true";
defparam \length[23] .power_up = "low";

dffeas \length[24] (
	.clk(outclk_wire_0),
	.d(in_data_reg_24),
	.asdata(\Add2~13_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[24]~q ),
	.prn(vcc));
defparam \length[24] .is_wysiwyg = "true";
defparam \length[24] .power_up = "low";

dffeas \length[25] (
	.clk(outclk_wire_0),
	.d(in_data_reg_25),
	.asdata(\Add2~17_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[25]~q ),
	.prn(vcc));
defparam \length[25] .is_wysiwyg = "true";
defparam \length[25] .power_up = "low";

dffeas \length[26] (
	.clk(outclk_wire_0),
	.d(in_data_reg_26),
	.asdata(\Add2~21_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[26]~q ),
	.prn(vcc));
defparam \length[26] .is_wysiwyg = "true";
defparam \length[26] .power_up = "low";

dffeas \length[12] (
	.clk(outclk_wire_0),
	.d(in_data_reg_12),
	.asdata(\Add2~25_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[12]~q ),
	.prn(vcc));
defparam \length[12] .is_wysiwyg = "true";
defparam \length[12] .power_up = "low";

dffeas \length[13] (
	.clk(outclk_wire_0),
	.d(in_data_reg_13),
	.asdata(\Add2~29_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[13]~q ),
	.prn(vcc));
defparam \length[13] .is_wysiwyg = "true";
defparam \length[13] .power_up = "low";

dffeas \length[14] (
	.clk(outclk_wire_0),
	.d(in_data_reg_14),
	.asdata(\Add2~33_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[14]~q ),
	.prn(vcc));
defparam \length[14] .is_wysiwyg = "true";
defparam \length[14] .power_up = "low";

dffeas \length[15] (
	.clk(outclk_wire_0),
	.d(in_data_reg_15),
	.asdata(\Add2~37_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[15]~q ),
	.prn(vcc));
defparam \length[15] .is_wysiwyg = "true";
defparam \length[15] .power_up = "low";

dffeas \length[16] (
	.clk(outclk_wire_0),
	.d(in_data_reg_16),
	.asdata(\Add2~41_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[16]~q ),
	.prn(vcc));
defparam \length[16] .is_wysiwyg = "true";
defparam \length[16] .power_up = "low";

dffeas \length[1] (
	.clk(outclk_wire_0),
	.d(in_data_reg_1),
	.asdata(\Add2~45_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[1]~q ),
	.prn(vcc));
defparam \length[1] .is_wysiwyg = "true";
defparam \length[1] .power_up = "low";

dffeas \length[2] (
	.clk(outclk_wire_0),
	.d(in_data_reg_2),
	.asdata(\Add2~49_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[2]~q ),
	.prn(vcc));
defparam \length[2] .is_wysiwyg = "true";
defparam \length[2] .power_up = "low";

dffeas \length[3] (
	.clk(outclk_wire_0),
	.d(in_data_reg_3),
	.asdata(\Add2~53_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[3]~q ),
	.prn(vcc));
defparam \length[3] .is_wysiwyg = "true";
defparam \length[3] .power_up = "low";

dffeas \length[4] (
	.clk(outclk_wire_0),
	.d(in_data_reg_4),
	.asdata(\Add2~57_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[4]~q ),
	.prn(vcc));
defparam \length[4] .is_wysiwyg = "true";
defparam \length[4] .power_up = "low";

dffeas \length[5] (
	.clk(outclk_wire_0),
	.d(in_data_reg_5),
	.asdata(\Add2~61_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[5]~q ),
	.prn(vcc));
defparam \length[5] .is_wysiwyg = "true";
defparam \length[5] .power_up = "low";

dffeas \length[6] (
	.clk(outclk_wire_0),
	.d(in_data_reg_6),
	.asdata(\Add2~65_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[6]~q ),
	.prn(vcc));
defparam \length[6] .is_wysiwyg = "true";
defparam \length[6] .power_up = "low";

dffeas \length[27] (
	.clk(outclk_wire_0),
	.d(in_data_reg_27),
	.asdata(\Add2~69_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[27]~q ),
	.prn(vcc));
defparam \length[27] .is_wysiwyg = "true";
defparam \length[27] .power_up = "low";

dffeas \length[28] (
	.clk(outclk_wire_0),
	.d(in_data_reg_28),
	.asdata(\Add2~73_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[28]~q ),
	.prn(vcc));
defparam \length[28] .is_wysiwyg = "true";
defparam \length[28] .power_up = "low";

dffeas \length[29] (
	.clk(outclk_wire_0),
	.d(in_data_reg_29),
	.asdata(\Add2~77_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[29]~q ),
	.prn(vcc));
defparam \length[29] .is_wysiwyg = "true";
defparam \length[29] .power_up = "low";

dffeas \length[11] (
	.clk(outclk_wire_0),
	.d(in_data_reg_11),
	.asdata(\Add2~81_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[11]~q ),
	.prn(vcc));
defparam \length[11] .is_wysiwyg = "true";
defparam \length[11] .power_up = "low";

dffeas \length[20] (
	.clk(outclk_wire_0),
	.d(in_data_reg_20),
	.asdata(\Add2~85_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[20]~q ),
	.prn(vcc));
defparam \length[20] .is_wysiwyg = "true";
defparam \length[20] .power_up = "low";

dffeas \length[21] (
	.clk(outclk_wire_0),
	.d(in_data_reg_21),
	.asdata(\Add2~89_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[21]~q ),
	.prn(vcc));
defparam \length[21] .is_wysiwyg = "true";
defparam \length[21] .power_up = "low";

dffeas \length[30] (
	.clk(outclk_wire_0),
	.d(in_data_reg_30),
	.asdata(\Add2~93_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[30]~q ),
	.prn(vcc));
defparam \length[30] .is_wysiwyg = "true";
defparam \length[30] .power_up = "low";

dffeas \length[17] (
	.clk(outclk_wire_0),
	.d(in_data_reg_17),
	.asdata(\Add2~97_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[17]~q ),
	.prn(vcc));
defparam \length[17] .is_wysiwyg = "true";
defparam \length[17] .power_up = "low";

dffeas \length[18] (
	.clk(outclk_wire_0),
	.d(in_data_reg_18),
	.asdata(\Add2~101_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[18]~q ),
	.prn(vcc));
defparam \length[18] .is_wysiwyg = "true";
defparam \length[18] .power_up = "low";

dffeas \length[19] (
	.clk(outclk_wire_0),
	.d(in_data_reg_19),
	.asdata(\Add2~105_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[19]~q ),
	.prn(vcc));
defparam \length[19] .is_wysiwyg = "true";
defparam \length[19] .power_up = "low";

dffeas \length[0] (
	.clk(outclk_wire_0),
	.d(in_data_reg_0),
	.asdata(\Add2~109_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[0]~q ),
	.prn(vcc));
defparam \length[0] .is_wysiwyg = "true";
defparam \length[0] .power_up = "low";

dffeas \length[7] (
	.clk(outclk_wire_0),
	.d(in_data_reg_7),
	.asdata(\Add2~113_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[7]~q ),
	.prn(vcc));
defparam \length[7] .is_wysiwyg = "true";
defparam \length[7] .power_up = "low";

dffeas \length[8] (
	.clk(outclk_wire_0),
	.d(in_data_reg_8),
	.asdata(\Add2~117_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[8]~q ),
	.prn(vcc));
defparam \length[8] .is_wysiwyg = "true";
defparam \length[8] .power_up = "low";

dffeas \length[9] (
	.clk(outclk_wire_0),
	.d(in_data_reg_9),
	.asdata(\Add2~121_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[9]~q ),
	.prn(vcc));
defparam \length[9] .is_wysiwyg = "true";
defparam \length[9] .power_up = "low";

dffeas \length[10] (
	.clk(outclk_wire_0),
	.d(in_data_reg_10),
	.asdata(\Add2~125_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\length[29]~0_combout ),
	.q(\length[10]~q ),
	.prn(vcc));
defparam \length[10] .is_wysiwyg = "true";
defparam \length[10] .power_up = "low";

cyclonev_lcell_comb \p1_writelength_eq_0~0 (
	.dataa(!\Add3~53_sumout ),
	.datab(!\Add3~57_sumout ),
	.datac(!\Add3~61_sumout ),
	.datad(!\Add3~65_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~0 .extended_lut = "off";
defparam \p1_writelength_eq_0~0 .lut_mask = 64'h8000800080008000;
defparam \p1_writelength_eq_0~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~1 (
	.dataa(!\Add3~33_sumout ),
	.datab(!\Add3~37_sumout ),
	.datac(!\Add3~41_sumout ),
	.datad(!\Add3~45_sumout ),
	.datae(!\Add3~49_sumout ),
	.dataf(!\p1_writelength_eq_0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~1 .extended_lut = "off";
defparam \p1_writelength_eq_0~1 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~2 (
	.dataa(!\Add3~13_sumout ),
	.datab(!\Add3~17_sumout ),
	.datac(!\Add3~21_sumout ),
	.datad(!\Add3~25_sumout ),
	.datae(!\Add3~29_sumout ),
	.dataf(!\p1_writelength_eq_0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~2 .extended_lut = "off";
defparam \p1_writelength_eq_0~2 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_done_write~0 (
	.dataa(!\writelength_eq_0~q ),
	.datab(!\Add3~1_sumout ),
	.datac(!\Add3~5_sumout ),
	.datad(!\Add3~9_sumout ),
	.datae(!\p1_writelength_eq_0~2_combout ),
	.dataf(!\p1_writelength_eq_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_done_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_done_write~0 .extended_lut = "off";
defparam \p1_done_write~0 .lut_mask = 64'hAAAAAAAAAAAAEAAA;
defparam \p1_done_write~0 .shared_arith = "off";

dffeas length_eq_0(
	.clk(outclk_wire_0),
	.d(\length_eq_0~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\length_eq_0~q ),
	.prn(vcc));
defparam length_eq_0.is_wysiwyg = "true";
defparam length_eq_0.power_up = "low";

cyclonev_lcell_comb \p1_length_eq_0~0 (
	.dataa(!\Add2~45_sumout ),
	.datab(!\Add2~49_sumout ),
	.datac(!\Add2~53_sumout ),
	.datad(!\Add2~57_sumout ),
	.datae(!\Add2~61_sumout ),
	.dataf(!\Add2~65_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~0 .extended_lut = "off";
defparam \p1_length_eq_0~0 .lut_mask = 64'h8000000000000000;
defparam \p1_length_eq_0~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~1 (
	.dataa(!\Add2~25_sumout ),
	.datab(!\Add2~29_sumout ),
	.datac(!\Add2~33_sumout ),
	.datad(!\Add2~37_sumout ),
	.datae(!\Add2~41_sumout ),
	.dataf(!\p1_length_eq_0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~1 .extended_lut = "off";
defparam \p1_length_eq_0~1 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~2 (
	.dataa(!\Add2~5_sumout ),
	.datab(!\Add2~9_sumout ),
	.datac(!\Add2~13_sumout ),
	.datad(!\Add2~17_sumout ),
	.datae(!\Add2~21_sumout ),
	.dataf(!\p1_length_eq_0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~2 .extended_lut = "off";
defparam \p1_length_eq_0~2 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~3 (
	.dataa(!\Add2~69_sumout ),
	.datab(!\Add2~73_sumout ),
	.datac(!\Add2~77_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~3 .extended_lut = "off";
defparam \p1_length_eq_0~3 .lut_mask = 64'h8080808080808080;
defparam \p1_length_eq_0~3 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~4 (
	.dataa(!\Add2~97_sumout ),
	.datab(!\Add2~101_sumout ),
	.datac(!\Add2~105_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~4 .extended_lut = "off";
defparam \p1_length_eq_0~4 .lut_mask = 64'h8080808080808080;
defparam \p1_length_eq_0~4 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~5 (
	.dataa(!f2h_ARREADY_0),
	.datab(!mem_used_7),
	.datac(!saved_grant_0),
	.datad(!WideOr1),
	.datae(!write),
	.dataf(!\length_eq_0~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~5 .extended_lut = "off";
defparam \p1_length_eq_0~5 .lut_mask = 64'h00000000000F0004;
defparam \p1_length_eq_0~5 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~6 (
	.dataa(!\Add2~109_sumout ),
	.datab(!\Add2~113_sumout ),
	.datac(!\Add2~117_sumout ),
	.datad(!\Add2~121_sumout ),
	.datae(!\Add2~125_sumout ),
	.dataf(!\p1_length_eq_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~6 .extended_lut = "off";
defparam \p1_length_eq_0~6 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~6 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~7 (
	.dataa(!\Add2~81_sumout ),
	.datab(!\Add2~85_sumout ),
	.datac(!\Add2~89_sumout ),
	.datad(!\Add2~93_sumout ),
	.datae(!\p1_length_eq_0~4_combout ),
	.dataf(!\p1_length_eq_0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~7 .extended_lut = "off";
defparam \p1_length_eq_0~7 .lut_mask = 64'h0000000000008000;
defparam \p1_length_eq_0~7 .shared_arith = "off";

cyclonev_lcell_comb \p1_done_read~0 (
	.dataa(!\length_eq_0~q ),
	.datab(!\Add2~1_sumout ),
	.datac(!\p1_length_eq_0~2_combout ),
	.datad(!\p1_length_eq_0~3_combout ),
	.datae(!\p1_length_eq_0~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_done_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_done_read~0 .extended_lut = "off";
defparam \p1_done_read~0 .lut_mask = 64'h5555555155555551;
defparam \p1_done_read~0 .shared_arith = "off";

cyclonev_lcell_comb \length_eq_0~0 (
	.dataa(!\length_eq_0~q ),
	.datab(!\Add2~1_sumout ),
	.datac(!\p1_length_eq_0~2_combout ),
	.datad(!\p1_length_eq_0~3_combout ),
	.datae(!\p1_length_eq_0~7_combout ),
	.dataf(!\p1_length~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\length_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \length_eq_0~0 .extended_lut = "off";
defparam \length_eq_0~0 .lut_mask = 64'hFFFFFFFF55555551;
defparam \length_eq_0~0 .shared_arith = "off";

cyclonev_lcell_comb \length[29]~0 (
	.dataa(!\p1_length_eq_0~5_combout ),
	.datab(!\p1_length~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\length[29]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \length[29]~0 .extended_lut = "off";
defparam \length[29]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \length[29]~0 .shared_arith = "off";

dffeas \readaddress[2] (
	.clk(outclk_wire_0),
	.d(\Add0~1_sumout ),
	.asdata(in_data_reg_2),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_2),
	.prn(vcc));
defparam \readaddress[2] .is_wysiwyg = "true";
defparam \readaddress[2] .power_up = "low";

dffeas \readaddress[3] (
	.clk(outclk_wire_0),
	.d(\Add0~5_sumout ),
	.asdata(in_data_reg_3),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_3),
	.prn(vcc));
defparam \readaddress[3] .is_wysiwyg = "true";
defparam \readaddress[3] .power_up = "low";

dffeas \readaddress[4] (
	.clk(outclk_wire_0),
	.d(\Add0~9_sumout ),
	.asdata(in_data_reg_4),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_4),
	.prn(vcc));
defparam \readaddress[4] .is_wysiwyg = "true";
defparam \readaddress[4] .power_up = "low";

dffeas \readaddress[5] (
	.clk(outclk_wire_0),
	.d(\Add0~13_sumout ),
	.asdata(in_data_reg_5),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_5),
	.prn(vcc));
defparam \readaddress[5] .is_wysiwyg = "true";
defparam \readaddress[5] .power_up = "low";

dffeas \readaddress[6] (
	.clk(outclk_wire_0),
	.d(\Add0~17_sumout ),
	.asdata(in_data_reg_6),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_6),
	.prn(vcc));
defparam \readaddress[6] .is_wysiwyg = "true";
defparam \readaddress[6] .power_up = "low";

dffeas \readaddress[7] (
	.clk(outclk_wire_0),
	.d(\Add0~21_sumout ),
	.asdata(in_data_reg_7),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_7),
	.prn(vcc));
defparam \readaddress[7] .is_wysiwyg = "true";
defparam \readaddress[7] .power_up = "low";

dffeas \readaddress[8] (
	.clk(outclk_wire_0),
	.d(\Add0~25_sumout ),
	.asdata(in_data_reg_8),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_8),
	.prn(vcc));
defparam \readaddress[8] .is_wysiwyg = "true";
defparam \readaddress[8] .power_up = "low";

dffeas \readaddress[9] (
	.clk(outclk_wire_0),
	.d(\Add0~29_sumout ),
	.asdata(in_data_reg_9),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_9),
	.prn(vcc));
defparam \readaddress[9] .is_wysiwyg = "true";
defparam \readaddress[9] .power_up = "low";

dffeas \readaddress[10] (
	.clk(outclk_wire_0),
	.d(\Add0~33_sumout ),
	.asdata(in_data_reg_10),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_10),
	.prn(vcc));
defparam \readaddress[10] .is_wysiwyg = "true";
defparam \readaddress[10] .power_up = "low";

dffeas \readaddress[11] (
	.clk(outclk_wire_0),
	.d(\Add0~37_sumout ),
	.asdata(in_data_reg_11),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_11),
	.prn(vcc));
defparam \readaddress[11] .is_wysiwyg = "true";
defparam \readaddress[11] .power_up = "low";

dffeas \readaddress[12] (
	.clk(outclk_wire_0),
	.d(\Add0~41_sumout ),
	.asdata(in_data_reg_12),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_12),
	.prn(vcc));
defparam \readaddress[12] .is_wysiwyg = "true";
defparam \readaddress[12] .power_up = "low";

dffeas \readaddress[13] (
	.clk(outclk_wire_0),
	.d(\Add0~45_sumout ),
	.asdata(in_data_reg_13),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_13),
	.prn(vcc));
defparam \readaddress[13] .is_wysiwyg = "true";
defparam \readaddress[13] .power_up = "low";

dffeas \readaddress[14] (
	.clk(outclk_wire_0),
	.d(\Add0~49_sumout ),
	.asdata(in_data_reg_14),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_14),
	.prn(vcc));
defparam \readaddress[14] .is_wysiwyg = "true";
defparam \readaddress[14] .power_up = "low";

dffeas \readaddress[15] (
	.clk(outclk_wire_0),
	.d(\Add0~53_sumout ),
	.asdata(in_data_reg_15),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_15),
	.prn(vcc));
defparam \readaddress[15] .is_wysiwyg = "true";
defparam \readaddress[15] .power_up = "low";

dffeas \readaddress[16] (
	.clk(outclk_wire_0),
	.d(\Add0~57_sumout ),
	.asdata(in_data_reg_16),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_16),
	.prn(vcc));
defparam \readaddress[16] .is_wysiwyg = "true";
defparam \readaddress[16] .power_up = "low";

dffeas \readaddress[17] (
	.clk(outclk_wire_0),
	.d(\Add0~61_sumout ),
	.asdata(in_data_reg_17),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_17),
	.prn(vcc));
defparam \readaddress[17] .is_wysiwyg = "true";
defparam \readaddress[17] .power_up = "low";

dffeas \readaddress[18] (
	.clk(outclk_wire_0),
	.d(\Add0~65_sumout ),
	.asdata(in_data_reg_18),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_18),
	.prn(vcc));
defparam \readaddress[18] .is_wysiwyg = "true";
defparam \readaddress[18] .power_up = "low";

dffeas \readaddress[19] (
	.clk(outclk_wire_0),
	.d(\Add0~69_sumout ),
	.asdata(in_data_reg_19),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_19),
	.prn(vcc));
defparam \readaddress[19] .is_wysiwyg = "true";
defparam \readaddress[19] .power_up = "low";

dffeas \readaddress[20] (
	.clk(outclk_wire_0),
	.d(\Add0~73_sumout ),
	.asdata(in_data_reg_20),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_20),
	.prn(vcc));
defparam \readaddress[20] .is_wysiwyg = "true";
defparam \readaddress[20] .power_up = "low";

dffeas \readaddress[21] (
	.clk(outclk_wire_0),
	.d(\Add0~77_sumout ),
	.asdata(in_data_reg_21),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_21),
	.prn(vcc));
defparam \readaddress[21] .is_wysiwyg = "true";
defparam \readaddress[21] .power_up = "low";

dffeas \readaddress[22] (
	.clk(outclk_wire_0),
	.d(\Add0~81_sumout ),
	.asdata(in_data_reg_22),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_22),
	.prn(vcc));
defparam \readaddress[22] .is_wysiwyg = "true";
defparam \readaddress[22] .power_up = "low";

dffeas \readaddress[23] (
	.clk(outclk_wire_0),
	.d(\Add0~85_sumout ),
	.asdata(in_data_reg_23),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_23),
	.prn(vcc));
defparam \readaddress[23] .is_wysiwyg = "true";
defparam \readaddress[23] .power_up = "low";

dffeas \readaddress[24] (
	.clk(outclk_wire_0),
	.d(\Add0~89_sumout ),
	.asdata(in_data_reg_24),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_24),
	.prn(vcc));
defparam \readaddress[24] .is_wysiwyg = "true";
defparam \readaddress[24] .power_up = "low";

dffeas \readaddress[25] (
	.clk(outclk_wire_0),
	.d(\Add0~93_sumout ),
	.asdata(in_data_reg_25),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_25),
	.prn(vcc));
defparam \readaddress[25] .is_wysiwyg = "true";
defparam \readaddress[25] .power_up = "low";

dffeas \readaddress[26] (
	.clk(outclk_wire_0),
	.d(\Add0~97_sumout ),
	.asdata(in_data_reg_26),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_26),
	.prn(vcc));
defparam \readaddress[26] .is_wysiwyg = "true";
defparam \readaddress[26] .power_up = "low";

dffeas \readaddress[27] (
	.clk(outclk_wire_0),
	.d(\Add0~101_sumout ),
	.asdata(in_data_reg_27),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_27),
	.prn(vcc));
defparam \readaddress[27] .is_wysiwyg = "true";
defparam \readaddress[27] .power_up = "low";

dffeas \readaddress[28] (
	.clk(outclk_wire_0),
	.d(\Add0~105_sumout ),
	.asdata(in_data_reg_28),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_28),
	.prn(vcc));
defparam \readaddress[28] .is_wysiwyg = "true";
defparam \readaddress[28] .power_up = "low";

dffeas \readaddress[29] (
	.clk(outclk_wire_0),
	.d(\Add0~109_sumout ),
	.asdata(in_data_reg_29),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_29),
	.prn(vcc));
defparam \readaddress[29] .is_wysiwyg = "true";
defparam \readaddress[29] .power_up = "low";

dffeas \readaddress[30] (
	.clk(outclk_wire_0),
	.d(\Add0~113_sumout ),
	.asdata(in_data_reg_30),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_30),
	.prn(vcc));
defparam \readaddress[30] .is_wysiwyg = "true";
defparam \readaddress[30] .power_up = "low";

dffeas \readaddress[31] (
	.clk(outclk_wire_0),
	.d(\Add0~117_sumout ),
	.asdata(in_data_reg_31),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(readaddress_31),
	.prn(vcc));
defparam \readaddress[31] .is_wysiwyg = "true";
defparam \readaddress[31] .power_up = "low";

dffeas \writeaddress[15] (
	.clk(outclk_wire_0),
	.d(\Add1~1_sumout ),
	.asdata(in_data_reg_15),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_15),
	.prn(vcc));
defparam \writeaddress[15] .is_wysiwyg = "true";
defparam \writeaddress[15] .power_up = "low";

dffeas \writeaddress[2] (
	.clk(outclk_wire_0),
	.d(\Add1~5_sumout ),
	.asdata(in_data_reg_2),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_2),
	.prn(vcc));
defparam \writeaddress[2] .is_wysiwyg = "true";
defparam \writeaddress[2] .power_up = "low";

dffeas \writeaddress[3] (
	.clk(outclk_wire_0),
	.d(\Add1~9_sumout ),
	.asdata(in_data_reg_3),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_3),
	.prn(vcc));
defparam \writeaddress[3] .is_wysiwyg = "true";
defparam \writeaddress[3] .power_up = "low";

dffeas \writeaddress[4] (
	.clk(outclk_wire_0),
	.d(\Add1~13_sumout ),
	.asdata(in_data_reg_4),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_4),
	.prn(vcc));
defparam \writeaddress[4] .is_wysiwyg = "true";
defparam \writeaddress[4] .power_up = "low";

dffeas \writeaddress[5] (
	.clk(outclk_wire_0),
	.d(\Add1~17_sumout ),
	.asdata(in_data_reg_5),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_5),
	.prn(vcc));
defparam \writeaddress[5] .is_wysiwyg = "true";
defparam \writeaddress[5] .power_up = "low";

dffeas \writeaddress[6] (
	.clk(outclk_wire_0),
	.d(\Add1~21_sumout ),
	.asdata(in_data_reg_6),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_6),
	.prn(vcc));
defparam \writeaddress[6] .is_wysiwyg = "true";
defparam \writeaddress[6] .power_up = "low";

dffeas \writeaddress[7] (
	.clk(outclk_wire_0),
	.d(\Add1~25_sumout ),
	.asdata(in_data_reg_7),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_7),
	.prn(vcc));
defparam \writeaddress[7] .is_wysiwyg = "true";
defparam \writeaddress[7] .power_up = "low";

dffeas \writeaddress[8] (
	.clk(outclk_wire_0),
	.d(\Add1~29_sumout ),
	.asdata(in_data_reg_8),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_8),
	.prn(vcc));
defparam \writeaddress[8] .is_wysiwyg = "true";
defparam \writeaddress[8] .power_up = "low";

dffeas \writeaddress[9] (
	.clk(outclk_wire_0),
	.d(\Add1~33_sumout ),
	.asdata(in_data_reg_9),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_9),
	.prn(vcc));
defparam \writeaddress[9] .is_wysiwyg = "true";
defparam \writeaddress[9] .power_up = "low";

dffeas \writeaddress[10] (
	.clk(outclk_wire_0),
	.d(\Add1~37_sumout ),
	.asdata(in_data_reg_10),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_10),
	.prn(vcc));
defparam \writeaddress[10] .is_wysiwyg = "true";
defparam \writeaddress[10] .power_up = "low";

dffeas \writeaddress[11] (
	.clk(outclk_wire_0),
	.d(\Add1~41_sumout ),
	.asdata(in_data_reg_11),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_11),
	.prn(vcc));
defparam \writeaddress[11] .is_wysiwyg = "true";
defparam \writeaddress[11] .power_up = "low";

dffeas \writeaddress[12] (
	.clk(outclk_wire_0),
	.d(\Add1~45_sumout ),
	.asdata(in_data_reg_12),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_12),
	.prn(vcc));
defparam \writeaddress[12] .is_wysiwyg = "true";
defparam \writeaddress[12] .power_up = "low";

dffeas \writeaddress[13] (
	.clk(outclk_wire_0),
	.d(\Add1~49_sumout ),
	.asdata(in_data_reg_13),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_13),
	.prn(vcc));
defparam \writeaddress[13] .is_wysiwyg = "true";
defparam \writeaddress[13] .power_up = "low";

dffeas \writeaddress[14] (
	.clk(outclk_wire_0),
	.d(\Add1~53_sumout ),
	.asdata(in_data_reg_14),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_14),
	.prn(vcc));
defparam \writeaddress[14] .is_wysiwyg = "true";
defparam \writeaddress[14] .power_up = "low";

dffeas \writeaddress[1] (
	.clk(outclk_wire_0),
	.d(\Add1~57_sumout ),
	.asdata(in_data_reg_1),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_1),
	.prn(vcc));
defparam \writeaddress[1] .is_wysiwyg = "true";
defparam \writeaddress[1] .power_up = "low";

dffeas \writeaddress[0] (
	.clk(outclk_wire_0),
	.d(\Add1~61_sumout ),
	.asdata(in_data_reg_0),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(writeaddress_0),
	.prn(vcc));
defparam \writeaddress[0] .is_wysiwyg = "true";
defparam \writeaddress[0] .power_up = "low";

dffeas \control[2] (
	.clk(outclk_wire_0),
	.d(\control[2]~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(control_2),
	.prn(vcc));
defparam \control[2] .is_wysiwyg = "true";
defparam \control[2] .power_up = "low";

dffeas \control[0] (
	.clk(outclk_wire_0),
	.d(in_data_reg_0),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(control_0),
	.prn(vcc));
defparam \control[0] .is_wysiwyg = "true";
defparam \control[0] .power_up = "low";

cyclonev_lcell_comb \write_writedata~0 (
	.dataa(!last_write_collision),
	.datab(!last_write_data_0),
	.datac(!q_b_0),
	.datad(!control_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~0 .extended_lut = "off";
defparam \write_writedata~0 .lut_mask = 64'h001B001B001B001B;
defparam \write_writedata~0 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~1 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_1),
	.datad(!q_b_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~1 .extended_lut = "off";
defparam \write_writedata~1 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~1 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~2 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_2),
	.datad(!q_b_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata2),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~2 .extended_lut = "off";
defparam \write_writedata~2 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~2 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~3 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_3),
	.datad(!q_b_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata3),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~3 .extended_lut = "off";
defparam \write_writedata~3 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~3 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~4 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_4),
	.datad(!q_b_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata4),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~4 .extended_lut = "off";
defparam \write_writedata~4 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~4 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~5 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_5),
	.datad(!q_b_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata5),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~5 .extended_lut = "off";
defparam \write_writedata~5 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~5 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~6 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_6),
	.datad(!q_b_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata6),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~6 .extended_lut = "off";
defparam \write_writedata~6 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~6 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~7 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_7),
	.datad(!q_b_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata7),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~7 .extended_lut = "off";
defparam \write_writedata~7 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~7 .shared_arith = "off";

dffeas \dma_ctl_readdata[0] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[0]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_0),
	.prn(vcc));
defparam \dma_ctl_readdata[0] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[0] .power_up = "low";

dffeas \dma_ctl_readdata[1] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[1]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_1),
	.prn(vcc));
defparam \dma_ctl_readdata[1] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[1] .power_up = "low";

dffeas \dma_ctl_readdata[2] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[2]~43_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_2),
	.prn(vcc));
defparam \dma_ctl_readdata[2] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[2] .power_up = "low";

dffeas \dma_ctl_readdata[3] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[3]~39_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_3),
	.prn(vcc));
defparam \dma_ctl_readdata[3] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[3] .power_up = "low";

dffeas \dma_ctl_readdata[4] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[4]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_4),
	.prn(vcc));
defparam \dma_ctl_readdata[4] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[4] .power_up = "low";

dffeas \dma_ctl_readdata[5] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[5]~35_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_5),
	.prn(vcc));
defparam \dma_ctl_readdata[5] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[5] .power_up = "low";

dffeas \dma_ctl_readdata[6] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[6]~31_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_6),
	.prn(vcc));
defparam \dma_ctl_readdata[6] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[6] .power_up = "low";

dffeas \dma_ctl_readdata[7] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[7]~27_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_7),
	.prn(vcc));
defparam \dma_ctl_readdata[7] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[7] .power_up = "low";

dffeas \dma_ctl_readdata[8] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[8]~23_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_8),
	.prn(vcc));
defparam \dma_ctl_readdata[8] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[8] .power_up = "low";

dffeas \dma_ctl_readdata[9] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[9]~19_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_9),
	.prn(vcc));
defparam \dma_ctl_readdata[9] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[9] .power_up = "low";

dffeas \dma_ctl_readdata[10] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[10]~15_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_10),
	.prn(vcc));
defparam \dma_ctl_readdata[10] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[10] .power_up = "low";

dffeas \dma_ctl_readdata[11] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[11]~11_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_11),
	.prn(vcc));
defparam \dma_ctl_readdata[11] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[11] .power_up = "low";

dffeas \dma_ctl_readdata[12] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[12]~7_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_12),
	.prn(vcc));
defparam \dma_ctl_readdata[12] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[12] .power_up = "low";

dffeas \dma_ctl_readdata[13] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[13]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_13),
	.prn(vcc));
defparam \dma_ctl_readdata[13] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[13] .power_up = "low";

dffeas \dma_ctl_readdata[14] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[14]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_14),
	.prn(vcc));
defparam \dma_ctl_readdata[14] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[14] .power_up = "low";

dffeas \dma_ctl_readdata[15] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[15]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_15),
	.prn(vcc));
defparam \dma_ctl_readdata[15] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[15] .power_up = "low";

dffeas \dma_ctl_readdata[16] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[16]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_16),
	.prn(vcc));
defparam \dma_ctl_readdata[16] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[16] .power_up = "low";

dffeas \dma_ctl_readdata[17] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[17]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_17),
	.prn(vcc));
defparam \dma_ctl_readdata[17] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[17] .power_up = "low";

dffeas \dma_ctl_readdata[18] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[18]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_18),
	.prn(vcc));
defparam \dma_ctl_readdata[18] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[18] .power_up = "low";

dffeas \dma_ctl_readdata[19] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[19]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_19),
	.prn(vcc));
defparam \dma_ctl_readdata[19] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[19] .power_up = "low";

dffeas \dma_ctl_readdata[20] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[20]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_20),
	.prn(vcc));
defparam \dma_ctl_readdata[20] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[20] .power_up = "low";

dffeas \dma_ctl_readdata[21] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[21]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_21),
	.prn(vcc));
defparam \dma_ctl_readdata[21] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[21] .power_up = "low";

dffeas \dma_ctl_readdata[22] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[22]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_22),
	.prn(vcc));
defparam \dma_ctl_readdata[22] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[22] .power_up = "low";

dffeas \dma_ctl_readdata[23] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[23]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_23),
	.prn(vcc));
defparam \dma_ctl_readdata[23] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[23] .power_up = "low";

dffeas \dma_ctl_readdata[24] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[24]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_24),
	.prn(vcc));
defparam \dma_ctl_readdata[24] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[24] .power_up = "low";

dffeas \dma_ctl_readdata[25] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[25]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_25),
	.prn(vcc));
defparam \dma_ctl_readdata[25] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[25] .power_up = "low";

dffeas \dma_ctl_readdata[26] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[26]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_26),
	.prn(vcc));
defparam \dma_ctl_readdata[26] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[26] .power_up = "low";

dffeas \dma_ctl_readdata[27] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[27]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_27),
	.prn(vcc));
defparam \dma_ctl_readdata[27] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[27] .power_up = "low";

dffeas \dma_ctl_readdata[28] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[28]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_28),
	.prn(vcc));
defparam \dma_ctl_readdata[28] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[28] .power_up = "low";

dffeas \dma_ctl_readdata[29] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[29]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_29),
	.prn(vcc));
defparam \dma_ctl_readdata[29] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[29] .power_up = "low";

dffeas \dma_ctl_readdata[30] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[30]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_30),
	.prn(vcc));
defparam \dma_ctl_readdata[30] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[30] .power_up = "low";

dffeas \dma_ctl_readdata[31] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[31]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_31),
	.prn(vcc));
defparam \dma_ctl_readdata[31] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[31] .power_up = "low";

cyclonev_lcell_comb \p1_readaddress~1 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_readaddress~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_readaddress~1 .extended_lut = "off";
defparam \p1_readaddress~1 .lut_mask = 64'h0008000800080008;
defparam \p1_readaddress~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~2 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~2 .extended_lut = "off";
defparam \Equal3~2 .lut_mask = 64'h1111111111111111;
defparam \Equal3~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_control~0 (
	.dataa(!\p1_readaddress~1_combout ),
	.datab(!\Equal3~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_control~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_control~0 .extended_lut = "off";
defparam \p1_control~0 .lut_mask = 64'h1111111111111111;
defparam \p1_control~0 .shared_arith = "off";

dffeas \control[12] (
	.clk(outclk_wire_0),
	.d(in_data_reg_12),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[12]~q ),
	.prn(vcc));
defparam \control[12] .is_wysiwyg = "true";
defparam \control[12] .power_up = "low";

cyclonev_lcell_comb \set_software_reset_bit~0 (
	.dataa(!\p1_readaddress~1_combout ),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!in_data_reg_12),
	.datad(!\Equal3~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\set_software_reset_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \set_software_reset_bit~0 .extended_lut = "off";
defparam \set_software_reset_bit~0 .lut_mask = 64'h0004000400040004;
defparam \set_software_reset_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \d1_softwarereset~0 (
	.dataa(!\software_reset_request~q ),
	.datab(!\control[12]~q ),
	.datac(!\d1_softwarereset~q ),
	.datad(!\set_software_reset_bit~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d1_softwarereset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d1_softwarereset~0 .extended_lut = "off";
defparam \d1_softwarereset~0 .lut_mask = 64'h0A220A220A220A22;
defparam \d1_softwarereset~0 .shared_arith = "off";

dffeas d1_softwarereset(
	.clk(outclk_wire_0),
	.d(\d1_softwarereset~0_combout ),
	.asdata(vcc),
	.clrn(!system_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d1_softwarereset~q ),
	.prn(vcc));
defparam d1_softwarereset.is_wysiwyg = "true";
defparam d1_softwarereset.power_up = "low";

cyclonev_lcell_comb \software_reset_request~0 (
	.dataa(!\software_reset_request~q ),
	.datab(!\d1_softwarereset~q ),
	.datac(!\set_software_reset_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\software_reset_request~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \software_reset_request~0 .extended_lut = "off";
defparam \software_reset_request~0 .lut_mask = 64'h0202020202020202;
defparam \software_reset_request~0 .shared_arith = "off";

dffeas software_reset_request(
	.clk(outclk_wire_0),
	.d(\software_reset_request~0_combout ),
	.asdata(vcc),
	.clrn(!system_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\software_reset_request~q ),
	.prn(vcc));
defparam software_reset_request.is_wysiwyg = "true";
defparam software_reset_request.power_up = "low";

cyclonev_lcell_comb \reset_n~0 (
	.dataa(!\software_reset_request~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reset_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reset_n~0 .extended_lut = "off";
defparam \reset_n~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reset_n~0 .shared_arith = "off";

dffeas reset_n(
	.clk(outclk_wire_0),
	.d(\reset_n~0_combout ),
	.asdata(vcc),
	.clrn(!system_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_n~q ),
	.prn(vcc));
defparam reset_n.is_wysiwyg = "true";
defparam reset_n.power_up = "low";

dffeas \control[8] (
	.clk(outclk_wire_0),
	.d(in_data_reg_8),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[8]~q ),
	.prn(vcc));
defparam \control[8] .is_wysiwyg = "true";
defparam \control[8] .power_up = "low";

cyclonev_lcell_comb \Add0~125 (
	.dataa(!control_0),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[8]~q ),
	.datae(gnd),
	.dataf(!\readaddress[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h0000FF0000005500;
defparam \Add0~125 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h4040404040404040;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_readaddress~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_readaddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_readaddress~0 .extended_lut = "off";
defparam \p1_readaddress~0 .lut_mask = 64'h0000000800000008;
defparam \p1_readaddress~0 .shared_arith = "off";

cyclonev_lcell_comb \readaddress[27]~0 (
	.dataa(!f2h_ARREADY_0),
	.datab(!mem_used_7),
	.datac(!saved_grant_0),
	.datad(!WideOr1),
	.datae(!write),
	.dataf(!\p1_readaddress~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readaddress[27]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readaddress[27]~0 .extended_lut = "off";
defparam \readaddress[27]~0 .lut_mask = 64'h000F0004FFFFFFFF;
defparam \readaddress[27]~0 .shared_arith = "off";

dffeas \readaddress[0] (
	.clk(outclk_wire_0),
	.d(\Add0~125_sumout ),
	.asdata(in_data_reg_0),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(\readaddress[0]~q ),
	.prn(vcc));
defparam \readaddress[0] .is_wysiwyg = "true";
defparam \readaddress[0] .power_up = "low";

cyclonev_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~121 .shared_arith = "off";

dffeas \readaddress[1] (
	.clk(outclk_wire_0),
	.d(\Add0~121_sumout ),
	.asdata(in_data_reg_1),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[27]~0_combout ),
	.q(\readaddress[1]~q ),
	.prn(vcc));
defparam \readaddress[1] .is_wysiwyg = "true";
defparam \readaddress[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!control_2),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[8]~q ),
	.datae(gnd),
	.dataf(!readaddress_2),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000AA00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~65 .shared_arith = "off";

cyclonev_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~69 .shared_arith = "off";

cyclonev_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~73 .shared_arith = "off";

cyclonev_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~77 .shared_arith = "off";

cyclonev_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~81 .shared_arith = "off";

cyclonev_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~85 .shared_arith = "off";

cyclonev_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~89 .shared_arith = "off";

cyclonev_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~93 .shared_arith = "off";

cyclonev_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~97 .shared_arith = "off";

cyclonev_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~101 .shared_arith = "off";

cyclonev_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~105 .shared_arith = "off";

cyclonev_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(\Add0~110 ),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~109 .shared_arith = "off";

cyclonev_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~113 .shared_arith = "off";

cyclonev_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~117 .shared_arith = "off";

dffeas \control[9] (
	.clk(outclk_wire_0),
	.d(in_data_reg_9),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[9]~q ),
	.prn(vcc));
defparam \control[9] .is_wysiwyg = "true";
defparam \control[9] .power_up = "low";

cyclonev_lcell_comb \Add1~61 (
	.dataa(!control_0),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[9]~q ),
	.datae(gnd),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~61_sumout ),
	.cout(\Add1~62 ),
	.shareout());
defparam \Add1~61 .extended_lut = "off";
defparam \Add1~61 .lut_mask = 64'h0000FF0000005500;
defparam \Add1~61 .shared_arith = "off";

cyclonev_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~57_sumout ),
	.cout(\Add1~58 ),
	.shareout());
defparam \Add1~57 .extended_lut = "off";
defparam \Add1~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~57 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!control_2),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[9]~q ),
	.datae(gnd),
	.dataf(!writeaddress_2),
	.datag(gnd),
	.cin(\Add1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF000000AA00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~37 .shared_arith = "off";

cyclonev_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout());
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~41 .shared_arith = "off";

cyclonev_lcell_comb \Add1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~45_sumout ),
	.cout(\Add1~46 ),
	.shareout());
defparam \Add1~45 .extended_lut = "off";
defparam \Add1~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~45 .shared_arith = "off";

cyclonev_lcell_comb \Add1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~49_sumout ),
	.cout(\Add1~50 ),
	.shareout());
defparam \Add1~49 .extended_lut = "off";
defparam \Add1~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~49 .shared_arith = "off";

cyclonev_lcell_comb \Add1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~53_sumout ),
	.cout(\Add1~54 ),
	.shareout());
defparam \Add1~53 .extended_lut = "off";
defparam \Add1~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~53 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~1 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~1 .extended_lut = "off";
defparam \Equal3~1 .lut_mask = 64'h0808080808080808;
defparam \Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_writeaddress~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writeaddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writeaddress~0 .extended_lut = "off";
defparam \p1_writeaddress~0 .lut_mask = 64'h0000000800000008;
defparam \p1_writeaddress~0 .shared_arith = "off";

cyclonev_lcell_comb \writeaddress[8]~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!wren),
	.datad(!in_data_reg_59),
	.datae(!mem),
	.dataf(!\Equal3~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writeaddress[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writeaddress[8]~0 .extended_lut = "off";
defparam \writeaddress[8]~0 .lut_mask = 64'h0F0F0F0F0F0F0F8F;
defparam \writeaddress[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \control[2]~0 (
	.dataa(!in_data_reg_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\control[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \control[2]~0 .extended_lut = "off";
defparam \control[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \control[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_0),
	.datad(!\writelength[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~109_sumout ),
	.cout(\Add3~110 ),
	.shareout(\Add3~111 ));
defparam \Add3~109 .extended_lut = "off";
defparam \Add3~109 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~109 .shared_arith = "on";

cyclonev_lcell_comb \Equal3~3 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~3 .extended_lut = "off";
defparam \Equal3~3 .lut_mask = 64'h0404040404040404;
defparam \Equal3~3 .shared_arith = "off";

cyclonev_lcell_comb \p1_length~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length~0 .extended_lut = "off";
defparam \p1_length~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \p1_length~0 .shared_arith = "off";

dffeas \writelength[30] (
	.clk(outclk_wire_0),
	.d(in_data_reg_30),
	.asdata(\Add3~5_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[30]~q ),
	.prn(vcc));
defparam \writelength[30] .is_wysiwyg = "true";
defparam \writelength[30] .power_up = "low";

cyclonev_lcell_comb \Add3~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~110 ),
	.sharein(\Add3~111 ),
	.combout(),
	.sumout(\Add3~113_sumout ),
	.cout(\Add3~114 ),
	.shareout(\Add3~115 ));
defparam \Add3~113 .extended_lut = "off";
defparam \Add3~113 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~113 .shared_arith = "on";

dffeas \writelength[1] (
	.clk(outclk_wire_0),
	.d(in_data_reg_1),
	.asdata(\Add3~113_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[1]~q ),
	.prn(vcc));
defparam \writelength[1] .is_wysiwyg = "true";
defparam \writelength[1] .power_up = "low";

cyclonev_lcell_comb \Add3~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_2),
	.datad(!\writelength[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~114 ),
	.sharein(\Add3~115 ),
	.combout(),
	.sumout(\Add3~117_sumout ),
	.cout(\Add3~118 ),
	.shareout(\Add3~119 ));
defparam \Add3~117 .extended_lut = "off";
defparam \Add3~117 .lut_mask = 64'h0000000F00000FF0;
defparam \Add3~117 .shared_arith = "on";

dffeas \writelength[2] (
	.clk(outclk_wire_0),
	.d(in_data_reg_2),
	.asdata(\Add3~117_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[2]~q ),
	.prn(vcc));
defparam \writelength[2] .is_wysiwyg = "true";
defparam \writelength[2] .power_up = "low";

cyclonev_lcell_comb \Add3~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~118 ),
	.sharein(\Add3~119 ),
	.combout(),
	.sumout(\Add3~121_sumout ),
	.cout(\Add3~122 ),
	.shareout(\Add3~123 ));
defparam \Add3~121 .extended_lut = "off";
defparam \Add3~121 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~121 .shared_arith = "on";

dffeas \writelength[3] (
	.clk(outclk_wire_0),
	.d(in_data_reg_3),
	.asdata(\Add3~121_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[3]~q ),
	.prn(vcc));
defparam \writelength[3] .is_wysiwyg = "true";
defparam \writelength[3] .power_up = "low";

cyclonev_lcell_comb \Add3~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~122 ),
	.sharein(\Add3~123 ),
	.combout(),
	.sumout(\Add3~125_sumout ),
	.cout(\Add3~126 ),
	.shareout(\Add3~127 ));
defparam \Add3~125 .extended_lut = "off";
defparam \Add3~125 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~125 .shared_arith = "on";

dffeas \writelength[4] (
	.clk(outclk_wire_0),
	.d(in_data_reg_4),
	.asdata(\Add3~125_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[4]~q ),
	.prn(vcc));
defparam \writelength[4] .is_wysiwyg = "true";
defparam \writelength[4] .power_up = "low";

cyclonev_lcell_comb \Add3~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~126 ),
	.sharein(\Add3~127 ),
	.combout(),
	.sumout(\Add3~53_sumout ),
	.cout(\Add3~54 ),
	.shareout(\Add3~55 ));
defparam \Add3~53 .extended_lut = "off";
defparam \Add3~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~53 .shared_arith = "on";

dffeas \writelength[5] (
	.clk(outclk_wire_0),
	.d(in_data_reg_5),
	.asdata(\Add3~53_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[5]~q ),
	.prn(vcc));
defparam \writelength[5] .is_wysiwyg = "true";
defparam \writelength[5] .power_up = "low";

cyclonev_lcell_comb \Add3~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~54 ),
	.sharein(\Add3~55 ),
	.combout(),
	.sumout(\Add3~57_sumout ),
	.cout(\Add3~58 ),
	.shareout(\Add3~59 ));
defparam \Add3~57 .extended_lut = "off";
defparam \Add3~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~57 .shared_arith = "on";

dffeas \writelength[6] (
	.clk(outclk_wire_0),
	.d(in_data_reg_6),
	.asdata(\Add3~57_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[6]~q ),
	.prn(vcc));
defparam \writelength[6] .is_wysiwyg = "true";
defparam \writelength[6] .power_up = "low";

cyclonev_lcell_comb \Add3~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~58 ),
	.sharein(\Add3~59 ),
	.combout(),
	.sumout(\Add3~61_sumout ),
	.cout(\Add3~62 ),
	.shareout(\Add3~63 ));
defparam \Add3~61 .extended_lut = "off";
defparam \Add3~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~61 .shared_arith = "on";

dffeas \writelength[7] (
	.clk(outclk_wire_0),
	.d(in_data_reg_7),
	.asdata(\Add3~61_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[7]~q ),
	.prn(vcc));
defparam \writelength[7] .is_wysiwyg = "true";
defparam \writelength[7] .power_up = "low";

cyclonev_lcell_comb \Add3~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~62 ),
	.sharein(\Add3~63 ),
	.combout(),
	.sumout(\Add3~65_sumout ),
	.cout(\Add3~66 ),
	.shareout(\Add3~67 ));
defparam \Add3~65 .extended_lut = "off";
defparam \Add3~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~65 .shared_arith = "on";

dffeas \writelength[8] (
	.clk(outclk_wire_0),
	.d(in_data_reg_8),
	.asdata(\Add3~65_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[8]~q ),
	.prn(vcc));
defparam \writelength[8] .is_wysiwyg = "true";
defparam \writelength[8] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~66 ),
	.sharein(\Add3~67 ),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout(\Add3~35 ));
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~33 .shared_arith = "on";

dffeas \writelength[9] (
	.clk(outclk_wire_0),
	.d(in_data_reg_9),
	.asdata(\Add3~33_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[9]~q ),
	.prn(vcc));
defparam \writelength[9] .is_wysiwyg = "true";
defparam \writelength[9] .power_up = "low";

cyclonev_lcell_comb \Add3~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(\Add3~35 ),
	.combout(),
	.sumout(\Add3~89_sumout ),
	.cout(\Add3~90 ),
	.shareout(\Add3~91 ));
defparam \Add3~89 .extended_lut = "off";
defparam \Add3~89 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~89 .shared_arith = "on";

dffeas \writelength[10] (
	.clk(outclk_wire_0),
	.d(in_data_reg_10),
	.asdata(\Add3~89_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[10]~q ),
	.prn(vcc));
defparam \writelength[10] .is_wysiwyg = "true";
defparam \writelength[10] .power_up = "low";

cyclonev_lcell_comb \Add3~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~90 ),
	.sharein(\Add3~91 ),
	.combout(),
	.sumout(\Add3~93_sumout ),
	.cout(\Add3~94 ),
	.shareout(\Add3~95 ));
defparam \Add3~93 .extended_lut = "off";
defparam \Add3~93 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~93 .shared_arith = "on";

dffeas \writelength[11] (
	.clk(outclk_wire_0),
	.d(in_data_reg_11),
	.asdata(\Add3~93_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[11]~q ),
	.prn(vcc));
defparam \writelength[11] .is_wysiwyg = "true";
defparam \writelength[11] .power_up = "low";

cyclonev_lcell_comb \Add3~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~94 ),
	.sharein(\Add3~95 ),
	.combout(),
	.sumout(\Add3~97_sumout ),
	.cout(\Add3~98 ),
	.shareout(\Add3~99 ));
defparam \Add3~97 .extended_lut = "off";
defparam \Add3~97 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~97 .shared_arith = "on";

dffeas \writelength[12] (
	.clk(outclk_wire_0),
	.d(in_data_reg_12),
	.asdata(\Add3~97_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[12]~q ),
	.prn(vcc));
defparam \writelength[12] .is_wysiwyg = "true";
defparam \writelength[12] .power_up = "low";

cyclonev_lcell_comb \Add3~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~98 ),
	.sharein(\Add3~99 ),
	.combout(),
	.sumout(\Add3~101_sumout ),
	.cout(\Add3~102 ),
	.shareout(\Add3~103 ));
defparam \Add3~101 .extended_lut = "off";
defparam \Add3~101 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~101 .shared_arith = "on";

dffeas \writelength[13] (
	.clk(outclk_wire_0),
	.d(in_data_reg_13),
	.asdata(\Add3~101_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[13]~q ),
	.prn(vcc));
defparam \writelength[13] .is_wysiwyg = "true";
defparam \writelength[13] .power_up = "low";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~102 ),
	.sharein(\Add3~103 ),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout(\Add3~39 ));
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~37 .shared_arith = "on";

dffeas \writelength[14] (
	.clk(outclk_wire_0),
	.d(in_data_reg_14),
	.asdata(\Add3~37_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[14]~q ),
	.prn(vcc));
defparam \writelength[14] .is_wysiwyg = "true";
defparam \writelength[14] .power_up = "low";

cyclonev_lcell_comb \Add3~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(\Add3~39 ),
	.combout(),
	.sumout(\Add3~105_sumout ),
	.cout(\Add3~106 ),
	.shareout(\Add3~107 ));
defparam \Add3~105 .extended_lut = "off";
defparam \Add3~105 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~105 .shared_arith = "on";

dffeas \writelength[15] (
	.clk(outclk_wire_0),
	.d(in_data_reg_15),
	.asdata(\Add3~105_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[15]~q ),
	.prn(vcc));
defparam \writelength[15] .is_wysiwyg = "true";
defparam \writelength[15] .power_up = "low";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~106 ),
	.sharein(\Add3~107 ),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout(\Add3~43 ));
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~41 .shared_arith = "on";

dffeas \writelength[16] (
	.clk(outclk_wire_0),
	.d(in_data_reg_16),
	.asdata(\Add3~41_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[16]~q ),
	.prn(vcc));
defparam \writelength[16] .is_wysiwyg = "true";
defparam \writelength[16] .power_up = "low";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(\Add3~43 ),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout(\Add3~47 ));
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~45 .shared_arith = "on";

dffeas \writelength[17] (
	.clk(outclk_wire_0),
	.d(in_data_reg_17),
	.asdata(\Add3~45_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[17]~q ),
	.prn(vcc));
defparam \writelength[17] .is_wysiwyg = "true";
defparam \writelength[17] .power_up = "low";

cyclonev_lcell_comb \Add3~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(\Add3~47 ),
	.combout(),
	.sumout(\Add3~49_sumout ),
	.cout(\Add3~50 ),
	.shareout(\Add3~51 ));
defparam \Add3~49 .extended_lut = "off";
defparam \Add3~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~49 .shared_arith = "on";

dffeas \writelength[18] (
	.clk(outclk_wire_0),
	.d(in_data_reg_18),
	.asdata(\Add3~49_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[18]~q ),
	.prn(vcc));
defparam \writelength[18] .is_wysiwyg = "true";
defparam \writelength[18] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~50 ),
	.sharein(\Add3~51 ),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout(\Add3~15 ));
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~13 .shared_arith = "on";

dffeas \writelength[19] (
	.clk(outclk_wire_0),
	.d(in_data_reg_19),
	.asdata(\Add3~13_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[19]~q ),
	.prn(vcc));
defparam \writelength[19] .is_wysiwyg = "true";
defparam \writelength[19] .power_up = "low";

cyclonev_lcell_comb \Add3~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(\Add3~15 ),
	.combout(),
	.sumout(\Add3~69_sumout ),
	.cout(\Add3~70 ),
	.shareout(\Add3~71 ));
defparam \Add3~69 .extended_lut = "off";
defparam \Add3~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~69 .shared_arith = "on";

dffeas \writelength[20] (
	.clk(outclk_wire_0),
	.d(in_data_reg_20),
	.asdata(\Add3~69_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[20]~q ),
	.prn(vcc));
defparam \writelength[20] .is_wysiwyg = "true";
defparam \writelength[20] .power_up = "low";

cyclonev_lcell_comb \Add3~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~70 ),
	.sharein(\Add3~71 ),
	.combout(),
	.sumout(\Add3~73_sumout ),
	.cout(\Add3~74 ),
	.shareout(\Add3~75 ));
defparam \Add3~73 .extended_lut = "off";
defparam \Add3~73 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~73 .shared_arith = "on";

dffeas \writelength[21] (
	.clk(outclk_wire_0),
	.d(in_data_reg_21),
	.asdata(\Add3~73_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[21]~q ),
	.prn(vcc));
defparam \writelength[21] .is_wysiwyg = "true";
defparam \writelength[21] .power_up = "low";

cyclonev_lcell_comb \Add3~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~74 ),
	.sharein(\Add3~75 ),
	.combout(),
	.sumout(\Add3~77_sumout ),
	.cout(\Add3~78 ),
	.shareout(\Add3~79 ));
defparam \Add3~77 .extended_lut = "off";
defparam \Add3~77 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~77 .shared_arith = "on";

dffeas \writelength[22] (
	.clk(outclk_wire_0),
	.d(in_data_reg_22),
	.asdata(\Add3~77_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[22]~q ),
	.prn(vcc));
defparam \writelength[22] .is_wysiwyg = "true";
defparam \writelength[22] .power_up = "low";

cyclonev_lcell_comb \Add3~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~78 ),
	.sharein(\Add3~79 ),
	.combout(),
	.sumout(\Add3~81_sumout ),
	.cout(\Add3~82 ),
	.shareout(\Add3~83 ));
defparam \Add3~81 .extended_lut = "off";
defparam \Add3~81 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~81 .shared_arith = "on";

dffeas \writelength[23] (
	.clk(outclk_wire_0),
	.d(in_data_reg_23),
	.asdata(\Add3~81_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[23]~q ),
	.prn(vcc));
defparam \writelength[23] .is_wysiwyg = "true";
defparam \writelength[23] .power_up = "low";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~82 ),
	.sharein(\Add3~83 ),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout(\Add3~19 ));
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~17 .shared_arith = "on";

dffeas \writelength[24] (
	.clk(outclk_wire_0),
	.d(in_data_reg_24),
	.asdata(\Add3~17_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[24]~q ),
	.prn(vcc));
defparam \writelength[24] .is_wysiwyg = "true";
defparam \writelength[24] .power_up = "low";

cyclonev_lcell_comb \Add3~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(\Add3~19 ),
	.combout(),
	.sumout(\Add3~85_sumout ),
	.cout(\Add3~86 ),
	.shareout(\Add3~87 ));
defparam \Add3~85 .extended_lut = "off";
defparam \Add3~85 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~85 .shared_arith = "on";

dffeas \writelength[25] (
	.clk(outclk_wire_0),
	.d(in_data_reg_25),
	.asdata(\Add3~85_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[25]~q ),
	.prn(vcc));
defparam \writelength[25] .is_wysiwyg = "true";
defparam \writelength[25] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~86 ),
	.sharein(\Add3~87 ),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout(\Add3~23 ));
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~21 .shared_arith = "on";

dffeas \writelength[26] (
	.clk(outclk_wire_0),
	.d(in_data_reg_26),
	.asdata(\Add3~21_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[26]~q ),
	.prn(vcc));
defparam \writelength[26] .is_wysiwyg = "true";
defparam \writelength[26] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(\Add3~23 ),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout(\Add3~27 ));
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~25 .shared_arith = "on";

dffeas \writelength[27] (
	.clk(outclk_wire_0),
	.d(in_data_reg_27),
	.asdata(\Add3~25_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[27]~q ),
	.prn(vcc));
defparam \writelength[27] .is_wysiwyg = "true";
defparam \writelength[27] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(\Add3~27 ),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout(\Add3~31 ));
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~29 .shared_arith = "on";

dffeas \writelength[28] (
	.clk(outclk_wire_0),
	.d(in_data_reg_28),
	.asdata(\Add3~29_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[28]~q ),
	.prn(vcc));
defparam \writelength[28] .is_wysiwyg = "true";
defparam \writelength[28] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(\Add3~31 ),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout(\Add3~3 ));
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~1 .shared_arith = "on";

dffeas \writelength[29] (
	.clk(outclk_wire_0),
	.d(in_data_reg_29),
	.asdata(\Add3~1_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[29]~q ),
	.prn(vcc));
defparam \writelength[29] .is_wysiwyg = "true";
defparam \writelength[29] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(\Add3~3 ),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout(\Add3~7 ));
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~5 .shared_arith = "on";

dffeas \writelength[31] (
	.clk(outclk_wire_0),
	.d(in_data_reg_31),
	.asdata(\Add3~9_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[31]~q ),
	.prn(vcc));
defparam \writelength[31] .is_wysiwyg = "true";
defparam \writelength[31] .power_up = "low";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(\Add3~7 ),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h000000000000FF00;
defparam \Add3~9 .shared_arith = "on";

cyclonev_lcell_comb \p1_writelength_eq_0~6 (
	.dataa(!\Add3~53_sumout ),
	.datab(!\Add3~57_sumout ),
	.datac(!\Add3~61_sumout ),
	.datad(!\Add3~65_sumout ),
	.datae(!\Add3~33_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~6 .extended_lut = "off";
defparam \p1_writelength_eq_0~6 .lut_mask = 64'h8000000080000000;
defparam \p1_writelength_eq_0~6 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~7 (
	.dataa(!\Add3~37_sumout ),
	.datab(!\Add3~41_sumout ),
	.datac(!\Add3~45_sumout ),
	.datad(!\Add3~49_sumout ),
	.datae(!\Add3~13_sumout ),
	.dataf(!\p1_writelength_eq_0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~7 .extended_lut = "off";
defparam \p1_writelength_eq_0~7 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~7 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~8 (
	.dataa(!\Add3~17_sumout ),
	.datab(!\Add3~21_sumout ),
	.datac(!\Add3~25_sumout ),
	.datad(!\Add3~29_sumout ),
	.datae(!\Add3~1_sumout ),
	.dataf(!\p1_writelength_eq_0~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~8 .extended_lut = "off";
defparam \p1_writelength_eq_0~8 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~8 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~3 (
	.dataa(!wren),
	.datab(!\Add3~109_sumout ),
	.datac(!\Add3~113_sumout ),
	.datad(!\Add3~117_sumout ),
	.datae(!\Add3~121_sumout ),
	.dataf(!\Add3~125_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~3 .extended_lut = "off";
defparam \p1_writelength_eq_0~3 .lut_mask = 64'h4000000000000000;
defparam \p1_writelength_eq_0~3 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~4 (
	.dataa(!\Add3~89_sumout ),
	.datab(!\Add3~93_sumout ),
	.datac(!\Add3~97_sumout ),
	.datad(!\Add3~101_sumout ),
	.datae(!\Add3~105_sumout ),
	.dataf(!\p1_writelength_eq_0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~4 .extended_lut = "off";
defparam \p1_writelength_eq_0~4 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~4 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~5 (
	.dataa(!\Add3~69_sumout ),
	.datab(!\Add3~73_sumout ),
	.datac(!\Add3~77_sumout ),
	.datad(!\Add3~81_sumout ),
	.datae(!\Add3~85_sumout ),
	.dataf(!\p1_writelength_eq_0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~5 .extended_lut = "off";
defparam \p1_writelength_eq_0~5 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~5 .shared_arith = "off";

cyclonev_lcell_comb \writelength_eq_0~0 (
	.dataa(!\writelength_eq_0~q ),
	.datab(!\Add3~5_sumout ),
	.datac(!\Add3~9_sumout ),
	.datad(!\p1_writelength_eq_0~8_combout ),
	.datae(!\p1_writelength_eq_0~5_combout ),
	.dataf(!\p1_length~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writelength_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writelength_eq_0~0 .extended_lut = "off";
defparam \writelength_eq_0~0 .lut_mask = 64'hFFFFFFFF55555515;
defparam \writelength_eq_0~0 .shared_arith = "off";

dffeas writelength_eq_0(
	.clk(outclk_wire_0),
	.d(\writelength_eq_0~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writelength_eq_0~q ),
	.prn(vcc));
defparam writelength_eq_0.is_wysiwyg = "true";
defparam writelength_eq_0.power_up = "low";

cyclonev_lcell_comb \writelength[13]~0 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_1),
	.datac(!mem_used_1),
	.datad(!fifo_empty),
	.datae(!\writelength_eq_0~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writelength[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writelength[13]~0 .extended_lut = "off";
defparam \writelength[13]~0 .lut_mask = 64'h0000001000000010;
defparam \writelength[13]~0 .shared_arith = "off";

cyclonev_lcell_comb \writelength[13]~1 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~3_combout ),
	.dataf(!\writelength[13]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writelength[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writelength[13]~1 .extended_lut = "off";
defparam \writelength[13]~1 .lut_mask = 64'h00000008FFFFFFFF;
defparam \writelength[13]~1 .shared_arith = "off";

dffeas \writelength[0] (
	.clk(outclk_wire_0),
	.d(in_data_reg_0),
	.asdata(\Add3~109_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_length~0_combout ),
	.ena(\writelength[13]~1_combout ),
	.q(\writelength[0]~q ),
	.prn(vcc));
defparam \writelength[0] .is_wysiwyg = "true";
defparam \writelength[0] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[0]~0 (
	.dataa(!writeaddress_0),
	.datab(!\readaddress[0]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[0]~0 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[0]~0 .lut_mask = 64'h0357035703570357;
defparam \p1_dma_ctl_readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~4 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!\Equal3~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~4 .extended_lut = "off";
defparam \Equal3~4 .lut_mask = 64'h2222222222222222;
defparam \Equal3~4 .shared_arith = "off";

dffeas \control[3] (
	.clk(outclk_wire_0),
	.d(in_data_reg_3),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[3]~q ),
	.prn(vcc));
defparam \control[3] .is_wysiwyg = "true";
defparam \control[3] .power_up = "low";

cyclonev_lcell_comb \control[7]~1 (
	.dataa(!in_data_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\control[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \control[7]~1 .extended_lut = "off";
defparam \control[7]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \control[7]~1 .shared_arith = "off";

dffeas \control[7] (
	.clk(outclk_wire_0),
	.d(\control[7]~1_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[7]~q ),
	.prn(vcc));
defparam \control[7] .is_wysiwyg = "true";
defparam \control[7] .power_up = "low";

cyclonev_lcell_comb \p1_done_write~1 (
	.dataa(!\control[7]~q ),
	.datab(!\writelength_eq_0~q ),
	.datac(!\Add3~5_sumout ),
	.datad(!\Add3~9_sumout ),
	.datae(!\p1_writelength_eq_0~8_combout ),
	.dataf(!\p1_writelength_eq_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_done_write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_done_write~1 .extended_lut = "off";
defparam \p1_done_write~1 .lut_mask = 64'h888888888888A888;
defparam \p1_done_write~1 .shared_arith = "off";

dffeas done_write(
	.clk(outclk_wire_0),
	.d(\p1_done_write~1_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\done_write~q ),
	.prn(vcc));
defparam done_write.is_wysiwyg = "true";
defparam done_write.power_up = "low";

cyclonev_lcell_comb done_transaction(
	.dataa(!\control[3]~q ),
	.datab(!\done_write~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\done_transaction~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam done_transaction.extended_lut = "off";
defparam done_transaction.lut_mask = 64'h1111111111111111;
defparam done_transaction.shared_arith = "off";

dffeas d1_done_transaction(
	.clk(outclk_wire_0),
	.d(\done_transaction~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d1_done_transaction~q ),
	.prn(vcc));
defparam d1_done_transaction.is_wysiwyg = "true";
defparam d1_done_transaction.power_up = "low";

cyclonev_lcell_comb flush_fifo(
	.dataa(!\control[3]~q ),
	.datab(!\done_write~q ),
	.datac(!\d1_done_transaction~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\flush_fifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam flush_fifo.extended_lut = "off";
defparam flush_fifo.lut_mask = 64'h1010101010101010;
defparam flush_fifo.shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata~1 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata~1 .extended_lut = "off";
defparam \p1_dma_ctl_readdata~1 .lut_mask = 64'h8080808080808080;
defparam \p1_dma_ctl_readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \done~0 (
	.dataa(!\flush_fifo~combout ),
	.datab(!\p1_readaddress~1_combout ),
	.datac(!\done~q ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \done~0 .extended_lut = "off";
defparam \done~0 .lut_mask = 64'h5F4C5F4C5F4C5F4C;
defparam \done~0 .shared_arith = "off";

dffeas done(
	.clk(outclk_wire_0),
	.d(\done~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\done~q ),
	.prn(vcc));
defparam done.is_wysiwyg = "true";
defparam done.power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[0]~2 (
	.dataa(!control_0),
	.datab(!\Equal3~4_combout ),
	.datac(!\done~q ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[0]~2 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[0]~2 .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[0] (
	.dataa(!\writelength[0]~q ),
	.datab(!\Equal3~3_combout ),
	.datac(!\p1_dma_ctl_readdata[0]~0_combout ),
	.datad(!\p1_dma_ctl_readdata[0]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[0] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[0] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \p1_dma_ctl_readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[1]~3 (
	.dataa(!writeaddress_1),
	.datab(!\readaddress[1]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[1]~3 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[1]~3 .lut_mask = 64'h0357035703570357;
defparam \p1_dma_ctl_readdata[1]~3 .shared_arith = "off";

dffeas \control[1] (
	.clk(outclk_wire_0),
	.d(in_data_reg_1),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[1]~q ),
	.prn(vcc));
defparam \control[1] .is_wysiwyg = "true";
defparam \control[1] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[1]~4 (
	.dataa(!\control[3]~q ),
	.datab(!\done_write~q ),
	.datac(!\Equal3~4_combout ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(!\control[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[1]~4 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[1]~4 .lut_mask = 64'h00440F4F00440F4F;
defparam \p1_dma_ctl_readdata[1]~4 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[1] (
	.dataa(!\writelength[1]~q ),
	.datab(!\Equal3~3_combout ),
	.datac(!\p1_dma_ctl_readdata[1]~3_combout ),
	.datad(!\p1_dma_ctl_readdata[1]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[1] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[1] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \p1_dma_ctl_readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[2]~43 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_2),
	.datad(!\writelength[2]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!control_2),
	.datag(!readaddress_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[2]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[2]~43 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[2]~43 .lut_mask = 64'h02024C6E0202082A;
defparam \p1_dma_ctl_readdata[2]~43 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[3]~39 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_3),
	.datad(!\writelength[3]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\control[3]~q ),
	.datag(!readaddress_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[3]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[3]~39 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[3]~39 .lut_mask = 64'h0202082A02024C6E;
defparam \p1_dma_ctl_readdata[3]~39 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[4]~5 (
	.dataa(!readaddress_4),
	.datab(!writeaddress_4),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[4]~5 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[4]~5 .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[4]~5 .shared_arith = "off";

dffeas \control[4] (
	.clk(outclk_wire_0),
	.d(in_data_reg_4),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[4]~q ),
	.prn(vcc));
defparam \control[4] .is_wysiwyg = "true";
defparam \control[4] .power_up = "low";

cyclonev_lcell_comb \len~0 (
	.dataa(!\writelength_eq_0~q ),
	.datab(!\flush_fifo~combout ),
	.datac(!\p1_readaddress~1_combout ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(!\len~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\len~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \len~0 .extended_lut = "off";
defparam \len~0 .lut_mask = 64'h2220FFF02220FFF0;
defparam \len~0 .shared_arith = "off";

dffeas len(
	.clk(outclk_wire_0),
	.d(\len~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\len~q ),
	.prn(vcc));
defparam len.is_wysiwyg = "true";
defparam len.power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[4]~6 (
	.dataa(!\Equal3~4_combout ),
	.datab(!\p1_dma_ctl_readdata~1_combout ),
	.datac(!\control[4]~q ),
	.datad(!\len~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[4]~6 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[4]~6 .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[4] (
	.dataa(!\writelength[4]~q ),
	.datab(!\Equal3~3_combout ),
	.datac(!\p1_dma_ctl_readdata[4]~5_combout ),
	.datad(!\p1_dma_ctl_readdata[4]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[4] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[4] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \p1_dma_ctl_readdata[4] .shared_arith = "off";

dffeas \control[5] (
	.clk(outclk_wire_0),
	.d(in_data_reg_5),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[5]~q ),
	.prn(vcc));
defparam \control[5] .is_wysiwyg = "true";
defparam \control[5] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[5]~35 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_5),
	.datad(!\control[5]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[5]~q ),
	.datag(!readaddress_5),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[5]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[5]~35 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[5]~35 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[5]~35 .shared_arith = "off";

dffeas \control[6] (
	.clk(outclk_wire_0),
	.d(in_data_reg_6),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[6]~q ),
	.prn(vcc));
defparam \control[6] .is_wysiwyg = "true";
defparam \control[6] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[6]~31 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_6),
	.datad(!\control[6]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[6]~q ),
	.datag(!readaddress_6),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[6]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[6]~31 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[6]~31 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[6]~31 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[7]~27 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_7),
	.datad(!\writelength[7]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\control[7]~q ),
	.datag(!readaddress_7),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[7]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[7]~27 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[7]~27 .lut_mask = 64'h02024C6E0202082A;
defparam \p1_dma_ctl_readdata[7]~27 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[8]~23 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_8),
	.datad(!\control[8]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[8]~q ),
	.datag(!readaddress_8),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[8]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[8]~23 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[8]~23 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[8]~23 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[9]~19 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_9),
	.datad(!\control[9]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[9]~q ),
	.datag(!readaddress_9),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[9]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[9]~19 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[9]~19 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[9]~19 .shared_arith = "off";

dffeas \control[10] (
	.clk(outclk_wire_0),
	.d(in_data_reg_10),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[10]~q ),
	.prn(vcc));
defparam \control[10] .is_wysiwyg = "true";
defparam \control[10] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[10]~15 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_10),
	.datad(!\control[10]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[10]~q ),
	.datag(!readaddress_10),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[10]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[10]~15 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[10]~15 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[10]~15 .shared_arith = "off";

dffeas \control[11] (
	.clk(outclk_wire_0),
	.d(in_data_reg_11),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[11]~q ),
	.prn(vcc));
defparam \control[11] .is_wysiwyg = "true";
defparam \control[11] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[11]~11 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_11),
	.datad(!\control[11]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[11]~q ),
	.datag(!readaddress_11),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[11]~11 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[11]~11 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[11]~11 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[12]~7 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_12),
	.datad(!\control[12]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[12]~q ),
	.datag(!readaddress_12),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[12]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[12]~7 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[12]~7 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[12]~7 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[13] (
	.dataa(!readaddress_13),
	.datab(!writeaddress_13),
	.datac(!\writelength[13]~q ),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(!int_nxt_addr_reg_dly_4),
	.dataf(!int_nxt_addr_reg_dly_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[13] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[13] .lut_mask = 64'h00550000330F0000;
defparam \p1_dma_ctl_readdata[13] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[14] (
	.dataa(!readaddress_14),
	.datab(!writeaddress_14),
	.datac(!\writelength[14]~q ),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(!int_nxt_addr_reg_dly_4),
	.dataf(!int_nxt_addr_reg_dly_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[14] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[14] .lut_mask = 64'h00550000330F0000;
defparam \p1_dma_ctl_readdata[14] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[15] (
	.dataa(!readaddress_15),
	.datab(!writeaddress_15),
	.datac(!\writelength[15]~q ),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(!int_nxt_addr_reg_dly_4),
	.dataf(!int_nxt_addr_reg_dly_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[15] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[15] .lut_mask = 64'h00550000330F0000;
defparam \p1_dma_ctl_readdata[15] .shared_arith = "off";

cyclonev_lcell_comb \Add1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~65_sumout ),
	.cout(\Add1~66 ),
	.shareout());
defparam \Add1~65 .extended_lut = "off";
defparam \Add1~65 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~65 .shared_arith = "off";

dffeas \writeaddress[16] (
	.clk(outclk_wire_0),
	.d(\Add1~65_sumout ),
	.asdata(in_data_reg_16),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[16]~q ),
	.prn(vcc));
defparam \writeaddress[16] .is_wysiwyg = "true";
defparam \writeaddress[16] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[16] (
	.dataa(!readaddress_16),
	.datab(!\writelength[16]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[16] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[16] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[16] .shared_arith = "off";

cyclonev_lcell_comb \Add1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~69_sumout ),
	.cout(\Add1~70 ),
	.shareout());
defparam \Add1~69 .extended_lut = "off";
defparam \Add1~69 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~69 .shared_arith = "off";

dffeas \writeaddress[17] (
	.clk(outclk_wire_0),
	.d(\Add1~69_sumout ),
	.asdata(in_data_reg_17),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[17]~q ),
	.prn(vcc));
defparam \writeaddress[17] .is_wysiwyg = "true";
defparam \writeaddress[17] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[17] (
	.dataa(!readaddress_17),
	.datab(!\writelength[17]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[17] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[17] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[17] .shared_arith = "off";

cyclonev_lcell_comb \Add1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~73_sumout ),
	.cout(\Add1~74 ),
	.shareout());
defparam \Add1~73 .extended_lut = "off";
defparam \Add1~73 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~73 .shared_arith = "off";

dffeas \writeaddress[18] (
	.clk(outclk_wire_0),
	.d(\Add1~73_sumout ),
	.asdata(in_data_reg_18),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[18]~q ),
	.prn(vcc));
defparam \writeaddress[18] .is_wysiwyg = "true";
defparam \writeaddress[18] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[18] (
	.dataa(!readaddress_18),
	.datab(!\writelength[18]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[18] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[18] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[18] .shared_arith = "off";

cyclonev_lcell_comb \Add1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~77_sumout ),
	.cout(\Add1~78 ),
	.shareout());
defparam \Add1~77 .extended_lut = "off";
defparam \Add1~77 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~77 .shared_arith = "off";

dffeas \writeaddress[19] (
	.clk(outclk_wire_0),
	.d(\Add1~77_sumout ),
	.asdata(in_data_reg_19),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[19]~q ),
	.prn(vcc));
defparam \writeaddress[19] .is_wysiwyg = "true";
defparam \writeaddress[19] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[19] (
	.dataa(!readaddress_19),
	.datab(!\writelength[19]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[19] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[19] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[19] .shared_arith = "off";

cyclonev_lcell_comb \Add1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~81_sumout ),
	.cout(\Add1~82 ),
	.shareout());
defparam \Add1~81 .extended_lut = "off";
defparam \Add1~81 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~81 .shared_arith = "off";

dffeas \writeaddress[20] (
	.clk(outclk_wire_0),
	.d(\Add1~81_sumout ),
	.asdata(in_data_reg_20),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[20]~q ),
	.prn(vcc));
defparam \writeaddress[20] .is_wysiwyg = "true";
defparam \writeaddress[20] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[20] (
	.dataa(!readaddress_20),
	.datab(!\writelength[20]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[20] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[20] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[20] .shared_arith = "off";

cyclonev_lcell_comb \Add1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~85_sumout ),
	.cout(\Add1~86 ),
	.shareout());
defparam \Add1~85 .extended_lut = "off";
defparam \Add1~85 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~85 .shared_arith = "off";

dffeas \writeaddress[21] (
	.clk(outclk_wire_0),
	.d(\Add1~85_sumout ),
	.asdata(in_data_reg_21),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[21]~q ),
	.prn(vcc));
defparam \writeaddress[21] .is_wysiwyg = "true";
defparam \writeaddress[21] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[21] (
	.dataa(!readaddress_21),
	.datab(!\writelength[21]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[21] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[21] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[21] .shared_arith = "off";

cyclonev_lcell_comb \Add1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~89_sumout ),
	.cout(\Add1~90 ),
	.shareout());
defparam \Add1~89 .extended_lut = "off";
defparam \Add1~89 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~89 .shared_arith = "off";

dffeas \writeaddress[22] (
	.clk(outclk_wire_0),
	.d(\Add1~89_sumout ),
	.asdata(in_data_reg_22),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[22]~q ),
	.prn(vcc));
defparam \writeaddress[22] .is_wysiwyg = "true";
defparam \writeaddress[22] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[22] (
	.dataa(!readaddress_22),
	.datab(!\writelength[22]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[22] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[22] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[22] .shared_arith = "off";

cyclonev_lcell_comb \Add1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~93_sumout ),
	.cout(\Add1~94 ),
	.shareout());
defparam \Add1~93 .extended_lut = "off";
defparam \Add1~93 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~93 .shared_arith = "off";

dffeas \writeaddress[23] (
	.clk(outclk_wire_0),
	.d(\Add1~93_sumout ),
	.asdata(in_data_reg_23),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[23]~q ),
	.prn(vcc));
defparam \writeaddress[23] .is_wysiwyg = "true";
defparam \writeaddress[23] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[23] (
	.dataa(!readaddress_23),
	.datab(!\writelength[23]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[23] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[23] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[23] .shared_arith = "off";

cyclonev_lcell_comb \Add1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~97_sumout ),
	.cout(\Add1~98 ),
	.shareout());
defparam \Add1~97 .extended_lut = "off";
defparam \Add1~97 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~97 .shared_arith = "off";

dffeas \writeaddress[24] (
	.clk(outclk_wire_0),
	.d(\Add1~97_sumout ),
	.asdata(in_data_reg_24),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[24]~q ),
	.prn(vcc));
defparam \writeaddress[24] .is_wysiwyg = "true";
defparam \writeaddress[24] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[24] (
	.dataa(!readaddress_24),
	.datab(!\writelength[24]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[24] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[24] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[24] .shared_arith = "off";

cyclonev_lcell_comb \Add1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~101_sumout ),
	.cout(\Add1~102 ),
	.shareout());
defparam \Add1~101 .extended_lut = "off";
defparam \Add1~101 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~101 .shared_arith = "off";

dffeas \writeaddress[25] (
	.clk(outclk_wire_0),
	.d(\Add1~101_sumout ),
	.asdata(in_data_reg_25),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[25]~q ),
	.prn(vcc));
defparam \writeaddress[25] .is_wysiwyg = "true";
defparam \writeaddress[25] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[25] (
	.dataa(!readaddress_25),
	.datab(!\writelength[25]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[25] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[25] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[25] .shared_arith = "off";

cyclonev_lcell_comb \Add1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~105_sumout ),
	.cout(\Add1~106 ),
	.shareout());
defparam \Add1~105 .extended_lut = "off";
defparam \Add1~105 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~105 .shared_arith = "off";

dffeas \writeaddress[26] (
	.clk(outclk_wire_0),
	.d(\Add1~105_sumout ),
	.asdata(in_data_reg_26),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[26]~q ),
	.prn(vcc));
defparam \writeaddress[26] .is_wysiwyg = "true";
defparam \writeaddress[26] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[26] (
	.dataa(!readaddress_26),
	.datab(!\writelength[26]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[26] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[26] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[26] .shared_arith = "off";

cyclonev_lcell_comb \Add1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writeaddress[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~109_sumout ),
	.cout(),
	.shareout());
defparam \Add1~109 .extended_lut = "off";
defparam \Add1~109 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~109 .shared_arith = "off";

dffeas \writeaddress[27] (
	.clk(outclk_wire_0),
	.d(\Add1~109_sumout ),
	.asdata(in_data_reg_27),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[8]~0_combout ),
	.q(\writeaddress[27]~q ),
	.prn(vcc));
defparam \writeaddress[27] .is_wysiwyg = "true";
defparam \writeaddress[27] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[27] (
	.dataa(!readaddress_27),
	.datab(!\writelength[27]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writeaddress[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[27] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[27] .lut_mask = 64'h050003000500F300;
defparam \p1_dma_ctl_readdata[27] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[28] (
	.dataa(!readaddress_28),
	.datab(!\writelength[28]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[28] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[28] .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[28] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[29] (
	.dataa(!readaddress_29),
	.datab(!\writelength[29]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[29] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[29] .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[29] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[30] (
	.dataa(!readaddress_30),
	.datab(!\writelength[30]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[30] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[30] .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[30] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[31] (
	.dataa(!readaddress_31),
	.datab(!\writelength[31]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[31] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[31] .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[31] .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_1_fifo_module (
	outclk_wire_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	fifo_empty1,
	wren,
	last_write_collision1,
	last_write_data_0,
	last_write_data_1,
	last_write_data_2,
	last_write_data_3,
	last_write_data_4,
	last_write_data_5,
	last_write_data_6,
	last_write_data_7,
	last_write_data_8,
	last_write_data_9,
	last_write_data_10,
	last_write_data_11,
	last_write_data_12,
	last_write_data_13,
	last_write_data_14,
	last_write_data_15,
	last_write_data_16,
	last_write_data_17,
	last_write_data_18,
	last_write_data_19,
	last_write_data_20,
	last_write_data_21,
	last_write_data_22,
	last_write_data_23,
	last_write_data_24,
	last_write_data_25,
	last_write_data_26,
	last_write_data_27,
	last_write_data_28,
	last_write_data_29,
	last_write_data_30,
	last_write_data_31,
	inc_read,
	flush_fifo,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	av_readdatavalid3,
	p1_fifo_full,
	reset_n,
	av_readdatavalid4,
	src0_valid,
	src_data_16,
	src_data_24,
	fifo_wr_data_0,
	src_data_17,
	src_data_25,
	fifo_wr_data_1,
	src_data_18,
	src_data_26,
	fifo_wr_data_2,
	src_data_19,
	src_data_27,
	fifo_wr_data_3,
	src_data_20,
	src_data_28,
	fifo_wr_data_4,
	src_data_21,
	src_data_29,
	fifo_wr_data_5,
	src_data_22,
	src_data_30,
	fifo_wr_data_6,
	src_data_23,
	src_data_31,
	fifo_wr_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	fifo_empty1;
input 	wren;
output 	last_write_collision1;
output 	last_write_data_0;
output 	last_write_data_1;
output 	last_write_data_2;
output 	last_write_data_3;
output 	last_write_data_4;
output 	last_write_data_5;
output 	last_write_data_6;
output 	last_write_data_7;
output 	last_write_data_8;
output 	last_write_data_9;
output 	last_write_data_10;
output 	last_write_data_11;
output 	last_write_data_12;
output 	last_write_data_13;
output 	last_write_data_14;
output 	last_write_data_15;
output 	last_write_data_16;
output 	last_write_data_17;
output 	last_write_data_18;
output 	last_write_data_19;
output 	last_write_data_20;
output 	last_write_data_21;
output 	last_write_data_22;
output 	last_write_data_23;
output 	last_write_data_24;
output 	last_write_data_25;
output 	last_write_data_26;
output 	last_write_data_27;
output 	last_write_data_28;
output 	last_write_data_29;
output 	last_write_data_30;
output 	last_write_data_31;
input 	inc_read;
input 	flush_fifo;
input 	av_readdatavalid;
input 	av_readdatavalid1;
input 	av_readdatavalid2;
input 	av_readdatavalid3;
output 	p1_fifo_full;
input 	reset_n;
input 	av_readdatavalid4;
input 	src0_valid;
input 	src_data_16;
input 	src_data_24;
input 	fifo_wr_data_0;
input 	src_data_17;
input 	src_data_25;
input 	fifo_wr_data_1;
input 	src_data_18;
input 	src_data_26;
input 	fifo_wr_data_2;
input 	src_data_19;
input 	src_data_27;
input 	fifo_wr_data_3;
input 	src_data_20;
input 	src_data_28;
input 	fifo_wr_data_4;
input 	src_data_21;
input 	src_data_29;
input 	fifo_wr_data_5;
input 	src_data_22;
input 	src_data_30;
input 	fifo_wr_data_6;
input 	src_data_23;
input 	src_data_31;
input 	fifo_wr_data_7;
input 	src_data_8;
input 	src_data_9;
input 	src_data_10;
input 	src_data_11;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rdaddress[0]~3_combout ;
wire \rdaddress_reg[0]~q ;
wire \rdaddress[1]~4_combout ;
wire \rdaddress_reg[1]~q ;
wire \rdaddress[2]~2_combout ;
wire \rdaddress_reg[2]~q ;
wire \Add1~0_combout ;
wire \rdaddress[3]~0_combout ;
wire \rdaddress_reg[3]~q ;
wire \Add1~1_combout ;
wire \rdaddress[4]~1_combout ;
wire \rdaddress_reg[4]~q ;
wire \wraddress~3_combout ;
wire \wraddress[3]~1_combout ;
wire \wraddress[0]~q ;
wire \wraddress~4_combout ;
wire \wraddress[1]~q ;
wire \wraddress~5_combout ;
wire \wraddress[2]~q ;
wire \wraddress~0_combout ;
wire \wraddress[3]~q ;
wire \wraddress~2_combout ;
wire \wraddress[4]~q ;
wire \p1_fifo_empty~0_combout ;
wire \p1_fifo_empty~1_combout ;
wire \p1_fifo_empty~2_combout ;
wire \p1_fifo_empty~3_combout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \write_collision~0_combout ;
wire \write_collision~combout ;
wire \last_write_collision~0_combout ;
wire \fifo_full~q ;
wire \estimated_wraddress~4_combout ;
wire \estimated_wraddress[4]~1_combout ;
wire \estimated_wraddress[0]~q ;
wire \estimated_wraddress~5_combout ;
wire \estimated_wraddress[1]~q ;
wire \estimated_wraddress~3_combout ;
wire \estimated_wraddress[2]~q ;
wire \estimated_wraddress~0_combout ;
wire \estimated_wraddress[3]~q ;
wire \estimated_wraddress~2_combout ;
wire \estimated_wraddress[4]~q ;
wire \p1_fifo_full~0_combout ;
wire \p1_fifo_full~1_combout ;
wire \p1_fifo_full~2_combout ;


Computer_System_Computer_System_dma_1_fifo_module_fifo_ram_module Computer_System_dma_1_fifo_module_fifo_ram(
	.outclk_wire_0(outclk_wire_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.av_readdatavalid(av_readdatavalid3),
	.rdaddress_3(\rdaddress[3]~0_combout ),
	.rdaddress_4(\rdaddress[4]~1_combout ),
	.rdaddress_2(\rdaddress[2]~2_combout ),
	.rdaddress_0(\rdaddress[0]~3_combout ),
	.rdaddress_1(\rdaddress[1]~4_combout ),
	.wraddress_3(\wraddress[3]~q ),
	.wraddress_4(\wraddress[4]~q ),
	.wraddress_0(\wraddress[0]~q ),
	.wraddress_1(\wraddress[1]~q ),
	.wraddress_2(\wraddress[2]~q ),
	.src_data_16(src_data_16),
	.src_data_24(src_data_24),
	.fifo_wr_data_0(fifo_wr_data_0),
	.src_data_17(src_data_17),
	.src_data_25(src_data_25),
	.fifo_wr_data_1(fifo_wr_data_1),
	.src_data_18(src_data_18),
	.src_data_26(src_data_26),
	.fifo_wr_data_2(fifo_wr_data_2),
	.src_data_19(src_data_19),
	.src_data_27(src_data_27),
	.fifo_wr_data_3(fifo_wr_data_3),
	.src_data_20(src_data_20),
	.src_data_28(src_data_28),
	.fifo_wr_data_4(fifo_wr_data_4),
	.src_data_21(src_data_21),
	.src_data_29(src_data_29),
	.fifo_wr_data_5(fifo_wr_data_5),
	.src_data_22(src_data_22),
	.src_data_30(src_data_30),
	.fifo_wr_data_6(fifo_wr_data_6),
	.src_data_23(src_data_23),
	.src_data_31(src_data_31),
	.fifo_wr_data_7(fifo_wr_data_7),
	.src_data_8(src_data_8),
	.src_data_9(src_data_9),
	.src_data_10(src_data_10),
	.src_data_11(src_data_11),
	.src_data_12(src_data_12),
	.src_data_13(src_data_13),
	.src_data_14(src_data_14),
	.src_data_15(src_data_15));

dffeas fifo_empty(
	.clk(outclk_wire_0),
	.d(\p1_fifo_empty~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_empty1),
	.prn(vcc));
defparam fifo_empty.is_wysiwyg = "true";
defparam fifo_empty.power_up = "low";

dffeas last_write_collision(
	.clk(outclk_wire_0),
	.d(\last_write_collision~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_write_collision1),
	.prn(vcc));
defparam last_write_collision.is_wysiwyg = "true";
defparam last_write_collision.power_up = "low";

dffeas \last_write_data[0] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_0),
	.prn(vcc));
defparam \last_write_data[0] .is_wysiwyg = "true";
defparam \last_write_data[0] .power_up = "low";

dffeas \last_write_data[1] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_1),
	.prn(vcc));
defparam \last_write_data[1] .is_wysiwyg = "true";
defparam \last_write_data[1] .power_up = "low";

dffeas \last_write_data[2] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_2),
	.prn(vcc));
defparam \last_write_data[2] .is_wysiwyg = "true";
defparam \last_write_data[2] .power_up = "low";

dffeas \last_write_data[3] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_3),
	.prn(vcc));
defparam \last_write_data[3] .is_wysiwyg = "true";
defparam \last_write_data[3] .power_up = "low";

dffeas \last_write_data[4] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_4),
	.prn(vcc));
defparam \last_write_data[4] .is_wysiwyg = "true";
defparam \last_write_data[4] .power_up = "low";

dffeas \last_write_data[5] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_5),
	.prn(vcc));
defparam \last_write_data[5] .is_wysiwyg = "true";
defparam \last_write_data[5] .power_up = "low";

dffeas \last_write_data[6] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_6),
	.prn(vcc));
defparam \last_write_data[6] .is_wysiwyg = "true";
defparam \last_write_data[6] .power_up = "low";

dffeas \last_write_data[7] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_7),
	.prn(vcc));
defparam \last_write_data[7] .is_wysiwyg = "true";
defparam \last_write_data[7] .power_up = "low";

dffeas \last_write_data[8] (
	.clk(outclk_wire_0),
	.d(src_data_8),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_8),
	.prn(vcc));
defparam \last_write_data[8] .is_wysiwyg = "true";
defparam \last_write_data[8] .power_up = "low";

dffeas \last_write_data[9] (
	.clk(outclk_wire_0),
	.d(src_data_9),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_9),
	.prn(vcc));
defparam \last_write_data[9] .is_wysiwyg = "true";
defparam \last_write_data[9] .power_up = "low";

dffeas \last_write_data[10] (
	.clk(outclk_wire_0),
	.d(src_data_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_10),
	.prn(vcc));
defparam \last_write_data[10] .is_wysiwyg = "true";
defparam \last_write_data[10] .power_up = "low";

dffeas \last_write_data[11] (
	.clk(outclk_wire_0),
	.d(src_data_11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_11),
	.prn(vcc));
defparam \last_write_data[11] .is_wysiwyg = "true";
defparam \last_write_data[11] .power_up = "low";

dffeas \last_write_data[12] (
	.clk(outclk_wire_0),
	.d(src_data_12),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_12),
	.prn(vcc));
defparam \last_write_data[12] .is_wysiwyg = "true";
defparam \last_write_data[12] .power_up = "low";

dffeas \last_write_data[13] (
	.clk(outclk_wire_0),
	.d(src_data_13),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_13),
	.prn(vcc));
defparam \last_write_data[13] .is_wysiwyg = "true";
defparam \last_write_data[13] .power_up = "low";

dffeas \last_write_data[14] (
	.clk(outclk_wire_0),
	.d(src_data_14),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_14),
	.prn(vcc));
defparam \last_write_data[14] .is_wysiwyg = "true";
defparam \last_write_data[14] .power_up = "low";

dffeas \last_write_data[15] (
	.clk(outclk_wire_0),
	.d(src_data_15),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_15),
	.prn(vcc));
defparam \last_write_data[15] .is_wysiwyg = "true";
defparam \last_write_data[15] .power_up = "low";

dffeas \last_write_data[16] (
	.clk(outclk_wire_0),
	.d(src_data_16),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_16),
	.prn(vcc));
defparam \last_write_data[16] .is_wysiwyg = "true";
defparam \last_write_data[16] .power_up = "low";

dffeas \last_write_data[17] (
	.clk(outclk_wire_0),
	.d(src_data_17),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_17),
	.prn(vcc));
defparam \last_write_data[17] .is_wysiwyg = "true";
defparam \last_write_data[17] .power_up = "low";

dffeas \last_write_data[18] (
	.clk(outclk_wire_0),
	.d(src_data_18),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_18),
	.prn(vcc));
defparam \last_write_data[18] .is_wysiwyg = "true";
defparam \last_write_data[18] .power_up = "low";

dffeas \last_write_data[19] (
	.clk(outclk_wire_0),
	.d(src_data_19),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_19),
	.prn(vcc));
defparam \last_write_data[19] .is_wysiwyg = "true";
defparam \last_write_data[19] .power_up = "low";

dffeas \last_write_data[20] (
	.clk(outclk_wire_0),
	.d(src_data_20),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_20),
	.prn(vcc));
defparam \last_write_data[20] .is_wysiwyg = "true";
defparam \last_write_data[20] .power_up = "low";

dffeas \last_write_data[21] (
	.clk(outclk_wire_0),
	.d(src_data_21),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_21),
	.prn(vcc));
defparam \last_write_data[21] .is_wysiwyg = "true";
defparam \last_write_data[21] .power_up = "low";

dffeas \last_write_data[22] (
	.clk(outclk_wire_0),
	.d(src_data_22),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_22),
	.prn(vcc));
defparam \last_write_data[22] .is_wysiwyg = "true";
defparam \last_write_data[22] .power_up = "low";

dffeas \last_write_data[23] (
	.clk(outclk_wire_0),
	.d(src_data_23),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_23),
	.prn(vcc));
defparam \last_write_data[23] .is_wysiwyg = "true";
defparam \last_write_data[23] .power_up = "low";

dffeas \last_write_data[24] (
	.clk(outclk_wire_0),
	.d(src_data_24),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_24),
	.prn(vcc));
defparam \last_write_data[24] .is_wysiwyg = "true";
defparam \last_write_data[24] .power_up = "low";

dffeas \last_write_data[25] (
	.clk(outclk_wire_0),
	.d(src_data_25),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_25),
	.prn(vcc));
defparam \last_write_data[25] .is_wysiwyg = "true";
defparam \last_write_data[25] .power_up = "low";

dffeas \last_write_data[26] (
	.clk(outclk_wire_0),
	.d(src_data_26),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_26),
	.prn(vcc));
defparam \last_write_data[26] .is_wysiwyg = "true";
defparam \last_write_data[26] .power_up = "low";

dffeas \last_write_data[27] (
	.clk(outclk_wire_0),
	.d(src_data_27),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_27),
	.prn(vcc));
defparam \last_write_data[27] .is_wysiwyg = "true";
defparam \last_write_data[27] .power_up = "low";

dffeas \last_write_data[28] (
	.clk(outclk_wire_0),
	.d(src_data_28),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_28),
	.prn(vcc));
defparam \last_write_data[28] .is_wysiwyg = "true";
defparam \last_write_data[28] .power_up = "low";

dffeas \last_write_data[29] (
	.clk(outclk_wire_0),
	.d(src_data_29),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_29),
	.prn(vcc));
defparam \last_write_data[29] .is_wysiwyg = "true";
defparam \last_write_data[29] .power_up = "low";

dffeas \last_write_data[30] (
	.clk(outclk_wire_0),
	.d(src_data_30),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_30),
	.prn(vcc));
defparam \last_write_data[30] .is_wysiwyg = "true";
defparam \last_write_data[30] .power_up = "low";

dffeas \last_write_data[31] (
	.clk(outclk_wire_0),
	.d(src_data_31),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_31),
	.prn(vcc));
defparam \last_write_data[31] .is_wysiwyg = "true";
defparam \last_write_data[31] .power_up = "low";

cyclonev_lcell_comb \p1_fifo_full~3 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\fifo_full~q ),
	.datad(!av_readdatavalid3),
	.datae(!\p1_fifo_full~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(p1_fifo_full),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~3 .extended_lut = "off";
defparam \p1_fifo_full~3 .lut_mask = 64'h080CCCCC080CCCCC;
defparam \p1_fifo_full~3 .shared_arith = "off";

cyclonev_lcell_comb \rdaddress[0]~3 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[0]~3 .extended_lut = "off";
defparam \rdaddress[0]~3 .lut_mask = 64'h4848484848484848;
defparam \rdaddress[0]~3 .shared_arith = "off";

dffeas \rdaddress_reg[0] (
	.clk(outclk_wire_0),
	.d(\rdaddress[0]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[0]~q ),
	.prn(vcc));
defparam \rdaddress_reg[0] .is_wysiwyg = "true";
defparam \rdaddress_reg[0] .power_up = "low";

cyclonev_lcell_comb \rdaddress[1]~4 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[0]~q ),
	.datad(!\rdaddress_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[1]~4 .extended_lut = "off";
defparam \rdaddress[1]~4 .lut_mask = 64'h408C408C408C408C;
defparam \rdaddress[1]~4 .shared_arith = "off";

dffeas \rdaddress_reg[1] (
	.clk(outclk_wire_0),
	.d(\rdaddress[1]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[1]~q ),
	.prn(vcc));
defparam \rdaddress_reg[1] .is_wysiwyg = "true";
defparam \rdaddress_reg[1] .power_up = "low";

cyclonev_lcell_comb \rdaddress[2]~2 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[0]~q ),
	.datad(!\rdaddress_reg[1]~q ),
	.datae(!\rdaddress_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[2]~2 .extended_lut = "off";
defparam \rdaddress[2]~2 .lut_mask = 64'h40008CCC40008CCC;
defparam \rdaddress[2]~2 .shared_arith = "off";

dffeas \rdaddress_reg[2] (
	.clk(outclk_wire_0),
	.d(\rdaddress[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[2]~q ),
	.prn(vcc));
defparam \rdaddress_reg[2] .is_wysiwyg = "true";
defparam \rdaddress_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\rdaddress_reg[0]~q ),
	.datab(!\rdaddress_reg[1]~q ),
	.datac(!\rdaddress_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8080808080808080;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \rdaddress[3]~0 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[3]~q ),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[3]~0 .extended_lut = "off";
defparam \rdaddress[3]~0 .lut_mask = 64'h0C480C480C480C48;
defparam \rdaddress[3]~0 .shared_arith = "off";

dffeas \rdaddress_reg[3] (
	.clk(outclk_wire_0),
	.d(\rdaddress[3]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[3]~q ),
	.prn(vcc));
defparam \rdaddress_reg[3] .is_wysiwyg = "true";
defparam \rdaddress_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\rdaddress_reg[0]~q ),
	.datab(!\rdaddress_reg[1]~q ),
	.datac(!\rdaddress_reg[2]~q ),
	.datad(!\rdaddress_reg[3]~q ),
	.datae(!\rdaddress_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h7FFF80007FFF8000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \rdaddress[4]~1 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[4]~q ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[4]~1 .extended_lut = "off";
defparam \rdaddress[4]~1 .lut_mask = 64'h4C084C084C084C08;
defparam \rdaddress[4]~1 .shared_arith = "off";

dffeas \rdaddress_reg[4] (
	.clk(outclk_wire_0),
	.d(\rdaddress[4]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[4]~q ),
	.prn(vcc));
defparam \rdaddress_reg[4] .is_wysiwyg = "true";
defparam \rdaddress_reg[4] .power_up = "low";

cyclonev_lcell_comb \wraddress~3 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~3 .extended_lut = "off";
defparam \wraddress~3 .lut_mask = 64'h8888888888888888;
defparam \wraddress~3 .shared_arith = "off";

cyclonev_lcell_comb \wraddress[3]~1 (
	.dataa(!src0_valid),
	.datab(!flush_fifo),
	.datac(!av_readdatavalid),
	.datad(!av_readdatavalid1),
	.datae(!av_readdatavalid2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress[3]~1 .extended_lut = "off";
defparam \wraddress[3]~1 .lut_mask = 64'h7773FFFF7773FFFF;
defparam \wraddress[3]~1 .shared_arith = "off";

dffeas \wraddress[0] (
	.clk(outclk_wire_0),
	.d(\wraddress~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[3]~1_combout ),
	.q(\wraddress[0]~q ),
	.prn(vcc));
defparam \wraddress[0] .is_wysiwyg = "true";
defparam \wraddress[0] .power_up = "low";

cyclonev_lcell_comb \wraddress~4 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~4 .extended_lut = "off";
defparam \wraddress~4 .lut_mask = 64'h8282828282828282;
defparam \wraddress~4 .shared_arith = "off";

dffeas \wraddress[1] (
	.clk(outclk_wire_0),
	.d(\wraddress~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[3]~1_combout ),
	.q(\wraddress[1]~q ),
	.prn(vcc));
defparam \wraddress[1] .is_wysiwyg = "true";
defparam \wraddress[1] .power_up = "low";

cyclonev_lcell_comb \wraddress~5 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\wraddress[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~5 .extended_lut = "off";
defparam \wraddress~5 .lut_mask = 64'h802A802A802A802A;
defparam \wraddress~5 .shared_arith = "off";

dffeas \wraddress[2] (
	.clk(outclk_wire_0),
	.d(\wraddress~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[3]~1_combout ),
	.q(\wraddress[2]~q ),
	.prn(vcc));
defparam \wraddress[2] .is_wysiwyg = "true";
defparam \wraddress[2] .power_up = "low";

cyclonev_lcell_comb \wraddress~0 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\wraddress[2]~q ),
	.datae(!\wraddress[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~0 .extended_lut = "off";
defparam \wraddress~0 .lut_mask = 64'h80002AAA80002AAA;
defparam \wraddress~0 .shared_arith = "off";

dffeas \wraddress[3] (
	.clk(outclk_wire_0),
	.d(\wraddress~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[3]~1_combout ),
	.q(\wraddress[3]~q ),
	.prn(vcc));
defparam \wraddress[3] .is_wysiwyg = "true";
defparam \wraddress[3] .power_up = "low";

cyclonev_lcell_comb \wraddress~2 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\wraddress[2]~q ),
	.datae(!\wraddress[3]~q ),
	.dataf(!\wraddress[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~2 .extended_lut = "off";
defparam \wraddress~2 .lut_mask = 64'h800000002AAAAAAA;
defparam \wraddress~2 .shared_arith = "off";

dffeas \wraddress[4] (
	.clk(outclk_wire_0),
	.d(\wraddress~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[3]~1_combout ),
	.q(\wraddress[4]~q ),
	.prn(vcc));
defparam \wraddress[4] .is_wysiwyg = "true";
defparam \wraddress[4] .power_up = "low";

cyclonev_lcell_comb \p1_fifo_empty~0 (
	.dataa(!\rdaddress_reg[0]~q ),
	.datab(!\rdaddress_reg[1]~q ),
	.datac(!\rdaddress_reg[2]~q ),
	.datad(!\wraddress[1]~q ),
	.datae(!\wraddress[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~0 .extended_lut = "off";
defparam \p1_fifo_empty~0 .lut_mask = 64'h6018068160180681;
defparam \p1_fifo_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_empty~1 (
	.dataa(!wren),
	.datab(!\rdaddress_reg[0]~q ),
	.datac(!\wraddress[0]~q ),
	.datad(!\p1_fifo_empty~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~1 .extended_lut = "off";
defparam \p1_fifo_empty~1 .lut_mask = 64'h0014001400140014;
defparam \p1_fifo_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_empty~2 (
	.dataa(!\rdaddress_reg[3]~q ),
	.datab(!\Add1~0_combout ),
	.datac(!\rdaddress_reg[4]~q ),
	.datad(!\wraddress[3]~q ),
	.datae(!\wraddress[4]~q ),
	.dataf(!\p1_fifo_empty~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~2 .extended_lut = "off";
defparam \p1_fifo_empty~2 .lut_mask = 64'h0000000090420924;
defparam \p1_fifo_empty~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_empty~3 (
	.dataa(!fifo_empty1),
	.datab(!flush_fifo),
	.datac(!av_readdatavalid3),
	.datad(!\p1_fifo_empty~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~3 .extended_lut = "off";
defparam \p1_fifo_empty~3 .lut_mask = 64'h4C0C4C0C4C0C4C0C;
defparam \p1_fifo_empty~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[0]~q ),
	.datad(!\rdaddress_reg[1]~q ),
	.datae(!\rdaddress_reg[2]~q ),
	.dataf(!\wraddress[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h40008CCCBFFF7333;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[3]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\wraddress[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h0C48F3B70C48F3B7;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~2 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[4]~q ),
	.datad(!\Add1~1_combout ),
	.datae(!\wraddress[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~2 .extended_lut = "off";
defparam \Equal2~2 .lut_mask = 64'h4C08B3F74C08B3F7;
defparam \Equal2~2 .shared_arith = "off";

cyclonev_lcell_comb \write_collision~0 (
	.dataa(!wren),
	.datab(!flush_fifo),
	.datac(!\rdaddress_reg[0]~q ),
	.datad(!\rdaddress_reg[1]~q ),
	.datae(!\wraddress[0]~q ),
	.dataf(!\wraddress[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_collision~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_collision~0 .extended_lut = "off";
defparam \write_collision~0 .lut_mask = 64'hB733084000844008;
defparam \write_collision~0 .shared_arith = "off";

cyclonev_lcell_comb write_collision(
	.dataa(!av_readdatavalid4),
	.datab(!av_readdatavalid2),
	.datac(!\Equal2~0_combout ),
	.datad(!\Equal2~1_combout ),
	.datae(!\Equal2~2_combout ),
	.dataf(!\write_collision~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_collision~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam write_collision.extended_lut = "off";
defparam write_collision.lut_mask = 64'h0000000070000000;
defparam write_collision.shared_arith = "off";

cyclonev_lcell_comb \last_write_collision~0 (
	.dataa(!wren),
	.datab(!last_write_collision1),
	.datac(!\write_collision~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_write_collision~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_write_collision~0 .extended_lut = "off";
defparam \last_write_collision~0 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \last_write_collision~0 .shared_arith = "off";

dffeas fifo_full(
	.clk(outclk_wire_0),
	.d(p1_fifo_full),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_full~q ),
	.prn(vcc));
defparam fifo_full.is_wysiwyg = "true";
defparam fifo_full.power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~4 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~4 .extended_lut = "off";
defparam \estimated_wraddress~4 .lut_mask = 64'h8888888888888888;
defparam \estimated_wraddress~4 .shared_arith = "off";

cyclonev_lcell_comb \estimated_wraddress[4]~1 (
	.dataa(!inc_read),
	.datab(!flush_fifo),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress[4]~1 .extended_lut = "off";
defparam \estimated_wraddress[4]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \estimated_wraddress[4]~1 .shared_arith = "off";

dffeas \estimated_wraddress[0] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[4]~1_combout ),
	.q(\estimated_wraddress[0]~q ),
	.prn(vcc));
defparam \estimated_wraddress[0] .is_wysiwyg = "true";
defparam \estimated_wraddress[0] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~5 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~5 .extended_lut = "off";
defparam \estimated_wraddress~5 .lut_mask = 64'h2828282828282828;
defparam \estimated_wraddress~5 .shared_arith = "off";

dffeas \estimated_wraddress[1] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[4]~1_combout ),
	.q(\estimated_wraddress[1]~q ),
	.prn(vcc));
defparam \estimated_wraddress[1] .is_wysiwyg = "true";
defparam \estimated_wraddress[1] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~3 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\estimated_wraddress[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~3 .extended_lut = "off";
defparam \estimated_wraddress~3 .lut_mask = 64'h02A802A802A802A8;
defparam \estimated_wraddress~3 .shared_arith = "off";

dffeas \estimated_wraddress[2] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[4]~1_combout ),
	.q(\estimated_wraddress[2]~q ),
	.prn(vcc));
defparam \estimated_wraddress[2] .is_wysiwyg = "true";
defparam \estimated_wraddress[2] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~0 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\estimated_wraddress[2]~q ),
	.datae(!\estimated_wraddress[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~0 .extended_lut = "off";
defparam \estimated_wraddress~0 .lut_mask = 64'h0002AAA80002AAA8;
defparam \estimated_wraddress~0 .shared_arith = "off";

dffeas \estimated_wraddress[3] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[4]~1_combout ),
	.q(\estimated_wraddress[3]~q ),
	.prn(vcc));
defparam \estimated_wraddress[3] .is_wysiwyg = "true";
defparam \estimated_wraddress[3] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~2 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\estimated_wraddress[2]~q ),
	.datae(!\estimated_wraddress[3]~q ),
	.dataf(!\estimated_wraddress[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~2 .extended_lut = "off";
defparam \estimated_wraddress~2 .lut_mask = 64'h00000002AAAAAAA8;
defparam \estimated_wraddress~2 .shared_arith = "off";

dffeas \estimated_wraddress[4] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[4]~1_combout ),
	.q(\estimated_wraddress[4]~q ),
	.prn(vcc));
defparam \estimated_wraddress[4] .is_wysiwyg = "true";
defparam \estimated_wraddress[4] .power_up = "low";

cyclonev_lcell_comb \p1_fifo_full~0 (
	.dataa(!\estimated_wraddress[0]~q ),
	.datab(!\rdaddress[0]~3_combout ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\rdaddress[1]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~0 .extended_lut = "off";
defparam \p1_fifo_full~0 .lut_mask = 64'h0660066006600660;
defparam \p1_fifo_full~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_full~1 (
	.dataa(!inc_read),
	.datab(!\estimated_wraddress[2]~q ),
	.datac(!\rdaddress[2]~2_combout ),
	.datad(!\p1_fifo_full~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~1 .extended_lut = "off";
defparam \p1_fifo_full~1 .lut_mask = 64'h0028002800280028;
defparam \p1_fifo_full~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_full~2 (
	.dataa(!\estimated_wraddress[3]~q ),
	.datab(!\rdaddress[3]~0_combout ),
	.datac(!\estimated_wraddress[4]~q ),
	.datad(!\rdaddress[4]~1_combout ),
	.datae(!\p1_fifo_full~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_full~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~2 .extended_lut = "off";
defparam \p1_fifo_full~2 .lut_mask = 64'h0000066000000660;
defparam \p1_fifo_full~2 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_1_fifo_module_fifo_ram_module (
	outclk_wire_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	av_readdatavalid,
	rdaddress_3,
	rdaddress_4,
	rdaddress_2,
	rdaddress_0,
	rdaddress_1,
	wraddress_3,
	wraddress_4,
	wraddress_0,
	wraddress_1,
	wraddress_2,
	src_data_16,
	src_data_24,
	fifo_wr_data_0,
	src_data_17,
	src_data_25,
	fifo_wr_data_1,
	src_data_18,
	src_data_26,
	fifo_wr_data_2,
	src_data_19,
	src_data_27,
	fifo_wr_data_3,
	src_data_20,
	src_data_28,
	fifo_wr_data_4,
	src_data_21,
	src_data_29,
	fifo_wr_data_5,
	src_data_22,
	src_data_30,
	fifo_wr_data_6,
	src_data_23,
	src_data_31,
	fifo_wr_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	av_readdatavalid;
input 	rdaddress_3;
input 	rdaddress_4;
input 	rdaddress_2;
input 	rdaddress_0;
input 	rdaddress_1;
input 	wraddress_3;
input 	wraddress_4;
input 	wraddress_0;
input 	wraddress_1;
input 	wraddress_2;
input 	src_data_16;
input 	src_data_24;
input 	fifo_wr_data_0;
input 	src_data_17;
input 	src_data_25;
input 	fifo_wr_data_1;
input 	src_data_18;
input 	src_data_26;
input 	fifo_wr_data_2;
input 	src_data_19;
input 	src_data_27;
input 	fifo_wr_data_3;
input 	src_data_20;
input 	src_data_28;
input 	fifo_wr_data_4;
input 	src_data_21;
input 	src_data_29;
input 	fifo_wr_data_5;
input 	src_data_22;
input 	src_data_30;
input 	fifo_wr_data_6;
input 	src_data_23;
input 	src_data_31;
input 	fifo_wr_data_7;
input 	src_data_8;
input 	src_data_9;
input 	src_data_10;
input 	src_data_11;
input 	src_data_12;
input 	src_data_13;
input 	src_data_14;
input 	src_data_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_lpm_ram_dp_1 lpm_ram_dp_component(
	.wrclock(outclk_wire_0),
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren(av_readdatavalid),
	.rdaddress({rdaddress_4,rdaddress_3,rdaddress_2,rdaddress_1,rdaddress_0}),
	.wraddress({wraddress_4,wraddress_3,wraddress_2,wraddress_1,wraddress_0}),
	.data({src_data_31,src_data_30,src_data_29,src_data_28,src_data_27,src_data_26,src_data_25,src_data_24,src_data_23,src_data_22,src_data_21,src_data_20,src_data_19,src_data_18,src_data_17,src_data_16,src_data_15,src_data_14,src_data_13,src_data_12,src_data_11,src_data_10,src_data_9,
src_data_8,fifo_wr_data_7,fifo_wr_data_6,fifo_wr_data_5,fifo_wr_data_4,fifo_wr_data_3,fifo_wr_data_2,fifo_wr_data_1,fifo_wr_data_0}));

endmodule

module Computer_System_lpm_ram_dp_1 (
	wrclock,
	q,
	wren,
	rdaddress,
	wraddress,
	data)/* synthesis synthesis_greybox=0 */;
input 	wrclock;
output 	[31:0] q;
input 	wren;
input 	[4:0] rdaddress;
input 	[4:0] wraddress;
input 	[31:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdpram_1 sram(
	.inclock(wrclock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren(wren),
	.rdaddress({rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.wraddress({wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module Computer_System_altdpram_1 (
	inclock,
	q,
	wren,
	rdaddress,
	wraddress,
	data)/* synthesis synthesis_greybox=0 */;
input 	inclock;
output 	[31:0] q;
input 	wren;
input 	[4:0] rdaddress;
input 	[4:0] wraddress;
input 	[31:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altsyncram_1 ram_block(
	.clock0(inclock),
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren_a(wren),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module Computer_System_altsyncram_1 (
	clock0,
	q_b,
	wren_a,
	address_b,
	address_a,
	data_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
output 	[31:0] q_b;
input 	wren_a;
input 	[13:0] address_b;
input 	[13:0] address_a;
input 	[31:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altsyncram_1j02 auto_generated(
	.clock0(clock0),
	.clock1(clock0),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}));

endmodule

module Computer_System_altsyncram_1j02 (
	clock0,
	clock1,
	q_b,
	wren_a,
	address_b,
	address_a,
	data_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
input 	clock1;
output 	[31:0] q_b;
input 	wren_a;
input 	[4:0] address_b;
input 	[4:0] address_a;
input 	[31:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.clk1_input_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.clk1_input_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.clk1_input_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.clk1_input_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.clk1_input_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.clk1_input_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.clk1_input_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.clk1_input_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.clk1_input_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.clk1_input_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.clk1_input_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.clk1_input_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.clk1_input_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.clk1_input_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.clk1_input_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.clk1_input_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Computer_System_dma_1:dma_1|Computer_System_dma_1_fifo_module:the_Computer_System_dma_1_fifo_module|Computer_System_dma_1_fifo_module_fifo_ram_module:Computer_System_dma_1_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module Computer_System_Computer_System_dma_1_mem_read (
	f2h_ARREADY_0,
	clk,
	mem_used_7,
	saved_grant_0,
	read_select1,
	hold_waitrequest,
	write,
	WideOr1,
	inc_read1,
	control_3,
	control_7,
	p1_done_write,
	p1_done_read,
	p1_fifo_full,
	reset_n)/* synthesis synthesis_greybox=0 */;
input 	f2h_ARREADY_0;
input 	clk;
input 	mem_used_7;
input 	saved_grant_0;
output 	read_select1;
input 	hold_waitrequest;
input 	write;
input 	WideOr1;
output 	inc_read1;
input 	control_3;
input 	control_7;
input 	p1_done_write;
input 	p1_done_read;
input 	p1_fifo_full;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Computer_System_dma_1_mem_read_idle~0_combout ;
wire \Computer_System_dma_1_mem_read_idle~4_combout ;
wire \Computer_System_dma_1_mem_read_idle~q ;
wire \Computer_System_dma_1_mem_read_access~0_combout ;
wire \p1_read_select~0_combout ;
wire \Computer_System_dma_1_mem_read_access~1_combout ;


dffeas read_select(
	.clk(clk),
	.d(\Computer_System_dma_1_mem_read_access~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_select1),
	.prn(vcc));
defparam read_select.is_wysiwyg = "true";
defparam read_select.power_up = "low";

cyclonev_lcell_comb inc_read(
	.dataa(!f2h_ARREADY_0),
	.datab(!mem_used_7),
	.datac(!saved_grant_0),
	.datad(!WideOr1),
	.datae(!write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(inc_read1),
	.sumout(),
	.cout(),
	.shareout());
defparam inc_read.extended_lut = "off";
defparam inc_read.lut_mask = 64'hFFF0FFFBFFF0FFFB;
defparam inc_read.shared_arith = "off";

cyclonev_lcell_comb \Computer_System_dma_1_mem_read_idle~0 (
	.dataa(!p1_fifo_full),
	.datab(!p1_done_read),
	.datac(!inc_read1),
	.datad(!p1_done_write),
	.datae(!\Computer_System_dma_1_mem_read_idle~q ),
	.dataf(!control_7),
	.datag(!control_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_1_mem_read_idle~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_1_mem_read_idle~0 .extended_lut = "on";
defparam \Computer_System_dma_1_mem_read_idle~0 .lut_mask = 64'hFDFFD0F0F5F55050;
defparam \Computer_System_dma_1_mem_read_idle~0 .shared_arith = "off";

cyclonev_lcell_comb \Computer_System_dma_1_mem_read_idle~4 (
	.dataa(!\Computer_System_dma_1_mem_read_idle~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_1_mem_read_idle~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_1_mem_read_idle~4 .extended_lut = "off";
defparam \Computer_System_dma_1_mem_read_idle~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Computer_System_dma_1_mem_read_idle~4 .shared_arith = "off";

dffeas Computer_System_dma_1_mem_read_idle(
	.clk(clk),
	.d(\Computer_System_dma_1_mem_read_idle~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\Computer_System_dma_1_mem_read_idle~q ),
	.prn(vcc));
defparam Computer_System_dma_1_mem_read_idle.is_wysiwyg = "true";
defparam Computer_System_dma_1_mem_read_idle.power_up = "low";

cyclonev_lcell_comb \Computer_System_dma_1_mem_read_access~0 (
	.dataa(!read_select1),
	.datab(!control_3),
	.datac(!\Computer_System_dma_1_mem_read_idle~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_1_mem_read_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_1_mem_read_access~0 .extended_lut = "off";
defparam \Computer_System_dma_1_mem_read_access~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \Computer_System_dma_1_mem_read_access~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_read_select~0 (
	.dataa(!f2h_ARREADY_0),
	.datab(!mem_used_7),
	.datac(!saved_grant_0),
	.datad(!read_select1),
	.datae(!hold_waitrequest),
	.dataf(!write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_read_select~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_read_select~0 .extended_lut = "off";
defparam \p1_read_select~0 .lut_mask = 64'h00FF00F000FF00FB;
defparam \p1_read_select~0 .shared_arith = "off";

cyclonev_lcell_comb \Computer_System_dma_1_mem_read_access~1 (
	.dataa(!\Computer_System_dma_1_mem_read_access~0_combout ),
	.datab(!control_7),
	.datac(!p1_done_write),
	.datad(!p1_done_read),
	.datae(!p1_fifo_full),
	.dataf(!\p1_read_select~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_1_mem_read_access~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_1_mem_read_access~1 .extended_lut = "off";
defparam \Computer_System_dma_1_mem_read_access~1 .lut_mask = 64'h22A20000FFFFFFFF;
defparam \Computer_System_dma_1_mem_read_access~1 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_1_read_data_mux (
	f2h_RVALID_0,
	clk,
	readaddress_0,
	readaddress_1,
	WideOr0,
	wait_latency_counter_1,
	control_2,
	control_0,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	reset_n,
	in_data_reg_59,
	mem,
	in_data_reg_3,
	src0_valid,
	src_data_8,
	src_data_81,
	src_data_16,
	src_data_24,
	src_data_0,
	src_data_01,
	fifo_wr_data_0,
	Equal3,
	src_data_9,
	src_data_91,
	src_data_17,
	src_data_25,
	src_data_1,
	src_data_11,
	fifo_wr_data_1,
	src_data_10,
	src_data_101,
	src_data_18,
	src_data_26,
	src_data_2,
	src_data_21,
	fifo_wr_data_2,
	src_data_111,
	src_data_112,
	src_data_19,
	src_data_27,
	src_data_3,
	src_data_31,
	fifo_wr_data_3,
	src_data_12,
	src_data_121,
	src_data_20,
	src_data_28,
	src_data_4,
	src_data_41,
	fifo_wr_data_4,
	src_data_13,
	src_data_131,
	src_data_211,
	src_data_29,
	src_data_5,
	src_data_51,
	fifo_wr_data_5,
	src_data_14,
	src_data_141,
	src_data_22,
	src_data_30,
	src_data_6,
	src_data_61,
	fifo_wr_data_6,
	src_data_15,
	src_data_151,
	src_data_23,
	src_data_311,
	src_data_7,
	src_data_71,
	fifo_wr_data_7,
	p1_length,
	control_8)/* synthesis synthesis_greybox=0 */;
input 	f2h_RVALID_0;
input 	clk;
input 	readaddress_0;
input 	readaddress_1;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	control_2;
input 	control_0;
input 	av_readdatavalid;
input 	av_readdatavalid1;
input 	av_readdatavalid2;
input 	reset_n;
input 	in_data_reg_59;
input 	mem;
input 	in_data_reg_3;
input 	src0_valid;
input 	src_data_8;
input 	src_data_81;
input 	src_data_16;
input 	src_data_24;
input 	src_data_0;
input 	src_data_01;
output 	fifo_wr_data_0;
input 	Equal3;
input 	src_data_9;
input 	src_data_91;
input 	src_data_17;
input 	src_data_25;
input 	src_data_1;
input 	src_data_11;
output 	fifo_wr_data_1;
input 	src_data_10;
input 	src_data_101;
input 	src_data_18;
input 	src_data_26;
input 	src_data_2;
input 	src_data_21;
output 	fifo_wr_data_2;
input 	src_data_111;
input 	src_data_112;
input 	src_data_19;
input 	src_data_27;
input 	src_data_3;
input 	src_data_31;
output 	fifo_wr_data_3;
input 	src_data_12;
input 	src_data_121;
input 	src_data_20;
input 	src_data_28;
input 	src_data_4;
input 	src_data_41;
output 	fifo_wr_data_4;
input 	src_data_13;
input 	src_data_131;
input 	src_data_211;
input 	src_data_29;
input 	src_data_5;
input 	src_data_51;
output 	fifo_wr_data_5;
input 	src_data_14;
input 	src_data_141;
input 	src_data_22;
input 	src_data_30;
input 	src_data_6;
input 	src_data_61;
output 	fifo_wr_data_6;
input 	src_data_15;
input 	src_data_151;
input 	src_data_23;
input 	src_data_311;
input 	src_data_7;
input 	src_data_71;
output 	fifo_wr_data_7;
input 	p1_length;
input 	control_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_data_mux_input~0_combout ;
wire \read_data_mux_input[0]~1_combout ;
wire \readdata_mux_select[1]~0_combout ;
wire \readdata_mux_select[0]~q ;
wire \Add0~0_combout ;
wire \read_data_mux_input[1]~2_combout ;
wire \readdata_mux_select[1]~q ;
wire \Equal4~0_combout ;
wire \fifo_wr_data~0_combout ;
wire \Equal4~1_combout ;
wire \fifo_wr_data[0]~1_combout ;
wire \fifo_wr_data[0]~2_combout ;
wire \fifo_wr_data~4_combout ;
wire \fifo_wr_data[1]~5_combout ;
wire \fifo_wr_data~7_combout ;
wire \fifo_wr_data[2]~8_combout ;
wire \fifo_wr_data~10_combout ;
wire \fifo_wr_data[3]~11_combout ;
wire \fifo_wr_data~13_combout ;
wire \fifo_wr_data[4]~14_combout ;
wire \fifo_wr_data~16_combout ;
wire \fifo_wr_data[5]~17_combout ;
wire \fifo_wr_data~19_combout ;
wire \fifo_wr_data[6]~20_combout ;
wire \fifo_wr_data~22_combout ;
wire \fifo_wr_data[7]~23_combout ;


cyclonev_lcell_comb \fifo_wr_data[0]~3 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\fifo_wr_data~0_combout ),
	.datac(!\Equal4~1_combout ),
	.datad(!src_data_16),
	.datae(!src_data_24),
	.dataf(!\fifo_wr_data[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[0]~3 .extended_lut = "off";
defparam \fifo_wr_data[0]~3 .lut_mask = 64'h333B373FFFFFFFFF;
defparam \fifo_wr_data[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[1]~6 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~4_combout ),
	.datad(!src_data_17),
	.datae(!src_data_25),
	.dataf(!\fifo_wr_data[1]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[1]~6 .extended_lut = "off";
defparam \fifo_wr_data[1]~6 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[2]~9 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~7_combout ),
	.datad(!src_data_18),
	.datae(!src_data_26),
	.dataf(!\fifo_wr_data[2]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[2]~9 .extended_lut = "off";
defparam \fifo_wr_data[2]~9 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[3]~12 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~10_combout ),
	.datad(!src_data_19),
	.datae(!src_data_27),
	.dataf(!\fifo_wr_data[3]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[3]~12 .extended_lut = "off";
defparam \fifo_wr_data[3]~12 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[3]~12 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[4]~15 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~13_combout ),
	.datad(!src_data_20),
	.datae(!src_data_28),
	.dataf(!\fifo_wr_data[4]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[4]~15 .extended_lut = "off";
defparam \fifo_wr_data[4]~15 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[4]~15 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[5]~18 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~16_combout ),
	.datad(!src_data_211),
	.datae(!src_data_29),
	.dataf(!\fifo_wr_data[5]~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[5]~18 .extended_lut = "off";
defparam \fifo_wr_data[5]~18 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[5]~18 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[6]~21 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~19_combout ),
	.datad(!src_data_22),
	.datae(!src_data_30),
	.dataf(!\fifo_wr_data[6]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[6]~21 .extended_lut = "off";
defparam \fifo_wr_data[6]~21 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[6]~21 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[7]~24 (
	.dataa(!\readdata_mux_select[0]~q ),
	.datab(!\Equal4~1_combout ),
	.datac(!\fifo_wr_data~22_combout ),
	.datad(!src_data_23),
	.datae(!src_data_311),
	.dataf(!\fifo_wr_data[7]~23_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[7]~24 .extended_lut = "off";
defparam \fifo_wr_data[7]~24 .lut_mask = 64'h0F2F1F3FFFFFFFFF;
defparam \fifo_wr_data[7]~24 .shared_arith = "off";

cyclonev_lcell_comb \read_data_mux_input~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!in_data_reg_3),
	.dataf(!Equal3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_data_mux_input~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_data_mux_input~0 .extended_lut = "off";
defparam \read_data_mux_input~0 .lut_mask = 64'h0000000000000008;
defparam \read_data_mux_input~0 .shared_arith = "off";

cyclonev_lcell_comb \read_data_mux_input[0]~1 (
	.dataa(!control_0),
	.datab(!control_8),
	.datac(!readaddress_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!p1_length),
	.dataf(!\read_data_mux_input~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_data_mux_input[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_data_mux_input[0]~1 .extended_lut = "off";
defparam \read_data_mux_input[0]~1 .lut_mask = 64'h0F0F44BB0F0F0F0F;
defparam \read_data_mux_input[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata_mux_select[1]~0 (
	.dataa(!src0_valid),
	.datab(!av_readdatavalid),
	.datac(!av_readdatavalid1),
	.datad(!av_readdatavalid2),
	.datae(!p1_length),
	.dataf(!\read_data_mux_input~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata_mux_select[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata_mux_select[1]~0 .extended_lut = "off";
defparam \readdata_mux_select[1]~0 .lut_mask = 64'hFFFF54FFFFFFFFFF;
defparam \readdata_mux_select[1]~0 .shared_arith = "off";

dffeas \readdata_mux_select[0] (
	.clk(clk),
	.d(\read_data_mux_input[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_mux_select[1]~0_combout ),
	.q(\readdata_mux_select[0]~q ),
	.prn(vcc));
defparam \readdata_mux_select[0] .is_wysiwyg = "true";
defparam \readdata_mux_select[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!control_0),
	.datab(!control_8),
	.datac(!\readdata_mux_select[0]~q ),
	.datad(!\readdata_mux_select[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h04FB04FB04FB04FB;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \read_data_mux_input[1]~2 (
	.dataa(!readaddress_1),
	.datab(!p1_length),
	.datac(!\read_data_mux_input~0_combout ),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_data_mux_input[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_data_mux_input[1]~2 .extended_lut = "off";
defparam \read_data_mux_input[1]~2 .lut_mask = 64'h4575457545754575;
defparam \read_data_mux_input[1]~2 .shared_arith = "off";

dffeas \readdata_mux_select[1] (
	.clk(clk),
	.d(\read_data_mux_input[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_mux_select[1]~0_combout ),
	.q(\readdata_mux_select[1]~q ),
	.prn(vcc));
defparam \readdata_mux_select[1] .is_wysiwyg = "true";
defparam \readdata_mux_select[1] .power_up = "low";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!control_0),
	.datab(!\readdata_mux_select[0]~q ),
	.datac(!\readdata_mux_select[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h1010101010101010;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_8),
	.datae(!src_data_81),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~0 .extended_lut = "off";
defparam \fifo_wr_data~0 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!control_0),
	.datab(!\readdata_mux_select[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h1111111111111111;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[0]~1 (
	.dataa(!control_2),
	.datab(!control_0),
	.datac(!\readdata_mux_select[0]~q ),
	.datad(!\readdata_mux_select[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[0]~1 .extended_lut = "off";
defparam \fifo_wr_data[0]~1 .lut_mask = 64'h4555455545554555;
defparam \fifo_wr_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[0]~2 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_0),
	.datae(!src_data_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[0]~2 .extended_lut = "off";
defparam \fifo_wr_data[0]~2 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~4 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_9),
	.datae(!src_data_91),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~4 .extended_lut = "off";
defparam \fifo_wr_data~4 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~4 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[1]~5 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_1),
	.datae(!src_data_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[1]~5 .extended_lut = "off";
defparam \fifo_wr_data[1]~5 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~7 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_10),
	.datae(!src_data_101),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~7 .extended_lut = "off";
defparam \fifo_wr_data~7 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~7 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[2]~8 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_2),
	.datae(!src_data_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[2]~8 .extended_lut = "off";
defparam \fifo_wr_data[2]~8 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[2]~8 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~10 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_111),
	.datae(!src_data_112),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~10 .extended_lut = "off";
defparam \fifo_wr_data~10 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~10 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[3]~11 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_3),
	.datae(!src_data_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[3]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[3]~11 .extended_lut = "off";
defparam \fifo_wr_data[3]~11 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[3]~11 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~13 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_12),
	.datae(!src_data_121),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~13 .extended_lut = "off";
defparam \fifo_wr_data~13 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~13 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[4]~14 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_4),
	.datae(!src_data_41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[4]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[4]~14 .extended_lut = "off";
defparam \fifo_wr_data[4]~14 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[4]~14 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~16 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_13),
	.datae(!src_data_131),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~16 .extended_lut = "off";
defparam \fifo_wr_data~16 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~16 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[5]~17 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_5),
	.datae(!src_data_51),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[5]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[5]~17 .extended_lut = "off";
defparam \fifo_wr_data[5]~17 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[5]~17 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~19 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_14),
	.datae(!src_data_141),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~19 .extended_lut = "off";
defparam \fifo_wr_data~19 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~19 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[6]~20 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_6),
	.datae(!src_data_61),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[6]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[6]~20 .extended_lut = "off";
defparam \fifo_wr_data[6]~20 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[6]~20 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~22 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\Equal4~0_combout ),
	.datad(!src_data_15),
	.datae(!src_data_151),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~22 .extended_lut = "off";
defparam \fifo_wr_data~22 .lut_mask = 64'h0003050700030507;
defparam \fifo_wr_data~22 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[7]~23 (
	.dataa(!f2h_RVALID_0),
	.datab(!src0_valid),
	.datac(!\fifo_wr_data[0]~1_combout ),
	.datad(!src_data_7),
	.datae(!src_data_71),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[7]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[7]~23 .extended_lut = "off";
defparam \fifo_wr_data[7]~23 .lut_mask = 64'h0030507000305070;
defparam \fifo_wr_data[7]~23 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_2 (
	f2h_AWREADY_0,
	f2h_WREADY_0,
	ram_block1a32,
	ram_block1a0,
	ram_block1a33,
	ram_block1a1,
	ram_block1a34,
	ram_block1a2,
	ram_block1a35,
	ram_block1a3,
	ram_block1a36,
	ram_block1a4,
	ram_block1a37,
	ram_block1a5,
	ram_block1a38,
	ram_block1a6,
	ram_block1a39,
	ram_block1a7,
	ram_block1a40,
	ram_block1a8,
	ram_block1a41,
	ram_block1a9,
	ram_block1a42,
	ram_block1a10,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a59,
	ram_block1a27,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	outclk_wire_0,
	writeaddress_2,
	writeaddress_3,
	writeaddress_4,
	writeaddress_5,
	writeaddress_6,
	writeaddress_7,
	writeaddress_8,
	writeaddress_9,
	writeaddress_10,
	writeaddress_11,
	writeaddress_12,
	writeaddress_13,
	writeaddress_14,
	writeaddress_15,
	writeaddress_16,
	writeaddress_17,
	writeaddress_18,
	writeaddress_19,
	writeaddress_20,
	writeaddress_21,
	writeaddress_22,
	writeaddress_23,
	writeaddress_24,
	writeaddress_25,
	writeaddress_26,
	writeaddress_27,
	writeaddress_28,
	writeaddress_29,
	writeaddress_30,
	writeaddress_31,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	writeaddress_1,
	writeaddress_0,
	readaddress_15,
	readaddress_2,
	readaddress_3,
	readaddress_4,
	readaddress_5,
	readaddress_6,
	readaddress_7,
	readaddress_8,
	readaddress_9,
	readaddress_10,
	readaddress_11,
	readaddress_12,
	readaddress_13,
	readaddress_14,
	hold_waitrequest,
	address_taken,
	mem_used_7,
	fifo_empty,
	src_valid,
	data_taken,
	last_write_collision,
	last_write_data_0,
	control_2,
	control_0,
	last_write_data_1,
	last_write_data_2,
	last_write_data_3,
	last_write_data_4,
	last_write_data_5,
	last_write_data_6,
	last_write_data_7,
	write_writedata,
	last_write_data_8,
	write_writedata1,
	last_write_data_9,
	write_writedata2,
	last_write_data_10,
	write_writedata3,
	last_write_data_11,
	write_writedata4,
	last_write_data_12,
	write_writedata5,
	last_write_data_13,
	write_writedata6,
	last_write_data_14,
	write_writedata7,
	last_write_data_15,
	last_write_data_16,
	last_write_data_17,
	last_write_data_18,
	last_write_data_19,
	last_write_data_20,
	last_write_data_21,
	last_write_data_22,
	last_write_data_23,
	last_write_data_24,
	last_write_data_25,
	last_write_data_26,
	last_write_data_27,
	last_write_data_28,
	last_write_data_29,
	last_write_data_30,
	last_write_data_31,
	WideOr0,
	wait_latency_counter_1,
	saved_grant_0,
	mem_used_1,
	system_reset_n,
	fifo_read,
	write_cp_ready,
	src0_valid,
	in_data_reg_2,
	in_data_reg_59,
	mem,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	address_reg_a_0,
	l1_w16_n0_mux_dataout,
	in_data_reg_0,
	l1_w17_n0_mux_dataout,
	l1_w18_n0_mux_dataout,
	l1_w19_n0_mux_dataout,
	l1_w20_n0_mux_dataout,
	l1_w21_n0_mux_dataout,
	l1_w22_n0_mux_dataout,
	l1_w23_n0_mux_dataout,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout,
	in_data_reg_1,
	dma_ctl_readdata_0,
	dma_ctl_readdata_1,
	dma_ctl_readdata_2,
	dma_ctl_readdata_3,
	dma_ctl_readdata_4,
	dma_ctl_readdata_5,
	dma_ctl_readdata_6,
	dma_ctl_readdata_7,
	dma_ctl_readdata_8,
	dma_ctl_readdata_9,
	dma_ctl_readdata_10,
	dma_ctl_readdata_11,
	dma_ctl_readdata_12,
	dma_ctl_readdata_13,
	dma_ctl_readdata_14,
	dma_ctl_readdata_15,
	dma_ctl_readdata_16,
	dma_ctl_readdata_17,
	dma_ctl_readdata_18,
	dma_ctl_readdata_19,
	dma_ctl_readdata_20,
	dma_ctl_readdata_21,
	dma_ctl_readdata_22,
	dma_ctl_readdata_23,
	dma_ctl_readdata_24,
	dma_ctl_readdata_25,
	dma_ctl_readdata_26,
	dma_ctl_readdata_27,
	dma_ctl_readdata_28,
	dma_ctl_readdata_29,
	dma_ctl_readdata_30,
	dma_ctl_readdata_31,
	read_select,
	read_latency_shift_reg)/* synthesis synthesis_greybox=0 */;
input 	f2h_AWREADY_0;
input 	f2h_WREADY_0;
input 	ram_block1a32;
input 	ram_block1a0;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a38;
input 	ram_block1a6;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a40;
input 	ram_block1a8;
input 	ram_block1a41;
input 	ram_block1a9;
input 	ram_block1a42;
input 	ram_block1a10;
input 	ram_block1a43;
input 	ram_block1a11;
input 	ram_block1a44;
input 	ram_block1a12;
input 	ram_block1a45;
input 	ram_block1a13;
input 	ram_block1a46;
input 	ram_block1a14;
input 	ram_block1a47;
input 	ram_block1a15;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	outclk_wire_0;
output 	writeaddress_2;
output 	writeaddress_3;
output 	writeaddress_4;
output 	writeaddress_5;
output 	writeaddress_6;
output 	writeaddress_7;
output 	writeaddress_8;
output 	writeaddress_9;
output 	writeaddress_10;
output 	writeaddress_11;
output 	writeaddress_12;
output 	writeaddress_13;
output 	writeaddress_14;
output 	writeaddress_15;
output 	writeaddress_16;
output 	writeaddress_17;
output 	writeaddress_18;
output 	writeaddress_19;
output 	writeaddress_20;
output 	writeaddress_21;
output 	writeaddress_22;
output 	writeaddress_23;
output 	writeaddress_24;
output 	writeaddress_25;
output 	writeaddress_26;
output 	writeaddress_27;
output 	writeaddress_28;
output 	writeaddress_29;
output 	writeaddress_30;
output 	writeaddress_31;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	writeaddress_1;
output 	writeaddress_0;
output 	readaddress_15;
output 	readaddress_2;
output 	readaddress_3;
output 	readaddress_4;
output 	readaddress_5;
output 	readaddress_6;
output 	readaddress_7;
output 	readaddress_8;
output 	readaddress_9;
output 	readaddress_10;
output 	readaddress_11;
output 	readaddress_12;
output 	readaddress_13;
output 	readaddress_14;
input 	hold_waitrequest;
input 	address_taken;
input 	mem_used_7;
output 	fifo_empty;
input 	src_valid;
input 	data_taken;
output 	last_write_collision;
output 	last_write_data_0;
output 	control_2;
output 	control_0;
output 	last_write_data_1;
output 	last_write_data_2;
output 	last_write_data_3;
output 	last_write_data_4;
output 	last_write_data_5;
output 	last_write_data_6;
output 	last_write_data_7;
output 	write_writedata;
output 	last_write_data_8;
output 	write_writedata1;
output 	last_write_data_9;
output 	write_writedata2;
output 	last_write_data_10;
output 	write_writedata3;
output 	last_write_data_11;
output 	write_writedata4;
output 	last_write_data_12;
output 	write_writedata5;
output 	last_write_data_13;
output 	write_writedata6;
output 	last_write_data_14;
output 	write_writedata7;
output 	last_write_data_15;
output 	last_write_data_16;
output 	last_write_data_17;
output 	last_write_data_18;
output 	last_write_data_19;
output 	last_write_data_20;
output 	last_write_data_21;
output 	last_write_data_22;
output 	last_write_data_23;
output 	last_write_data_24;
output 	last_write_data_25;
output 	last_write_data_26;
output 	last_write_data_27;
output 	last_write_data_28;
output 	last_write_data_29;
output 	last_write_data_30;
output 	last_write_data_31;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	saved_grant_0;
input 	mem_used_1;
input 	system_reset_n;
output 	fifo_read;
input 	write_cp_ready;
input 	src0_valid;
input 	in_data_reg_2;
input 	in_data_reg_59;
input 	mem;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_4;
input 	int_nxt_addr_reg_dly_3;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
input 	address_reg_a_0;
input 	l1_w16_n0_mux_dataout;
input 	in_data_reg_0;
input 	l1_w17_n0_mux_dataout;
input 	l1_w18_n0_mux_dataout;
input 	l1_w19_n0_mux_dataout;
input 	l1_w20_n0_mux_dataout;
input 	l1_w21_n0_mux_dataout;
input 	l1_w22_n0_mux_dataout;
input 	l1_w23_n0_mux_dataout;
input 	l1_w8_n0_mux_dataout;
input 	l1_w9_n0_mux_dataout;
input 	l1_w10_n0_mux_dataout;
input 	l1_w11_n0_mux_dataout;
input 	l1_w12_n0_mux_dataout;
input 	l1_w13_n0_mux_dataout;
input 	l1_w14_n0_mux_dataout;
input 	l1_w15_n0_mux_dataout;
input 	l1_w24_n0_mux_dataout;
input 	l1_w25_n0_mux_dataout;
input 	l1_w26_n0_mux_dataout;
input 	l1_w27_n0_mux_dataout;
input 	l1_w28_n0_mux_dataout;
input 	l1_w29_n0_mux_dataout;
input 	l1_w30_n0_mux_dataout;
input 	l1_w31_n0_mux_dataout;
input 	in_data_reg_1;
output 	dma_ctl_readdata_0;
output 	dma_ctl_readdata_1;
output 	dma_ctl_readdata_2;
output 	dma_ctl_readdata_3;
output 	dma_ctl_readdata_4;
output 	dma_ctl_readdata_5;
output 	dma_ctl_readdata_6;
output 	dma_ctl_readdata_7;
output 	dma_ctl_readdata_8;
output 	dma_ctl_readdata_9;
output 	dma_ctl_readdata_10;
output 	dma_ctl_readdata_11;
output 	dma_ctl_readdata_12;
output 	dma_ctl_readdata_13;
output 	dma_ctl_readdata_14;
output 	dma_ctl_readdata_15;
output 	dma_ctl_readdata_16;
output 	dma_ctl_readdata_17;
output 	dma_ctl_readdata_18;
output 	dma_ctl_readdata_19;
output 	dma_ctl_readdata_20;
output 	dma_ctl_readdata_21;
output 	dma_ctl_readdata_22;
output 	dma_ctl_readdata_23;
output 	dma_ctl_readdata_24;
output 	dma_ctl_readdata_25;
output 	dma_ctl_readdata_26;
output 	dma_ctl_readdata_27;
output 	dma_ctl_readdata_28;
output 	dma_ctl_readdata_29;
output 	dma_ctl_readdata_30;
output 	dma_ctl_readdata_31;
output 	read_select;
input 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add2~1_sumout ;
wire \Add2~2 ;
wire \Add2~3 ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add2~7 ;
wire \Add2~9_sumout ;
wire \Add2~13_sumout ;
wire \Add2~14 ;
wire \Add2~15 ;
wire \Add2~17_sumout ;
wire \Add2~18 ;
wire \Add2~19 ;
wire \Add2~21_sumout ;
wire \Add2~22 ;
wire \Add2~23 ;
wire \Add2~25_sumout ;
wire \Add2~26 ;
wire \Add2~27 ;
wire \Add2~29_sumout ;
wire \Add2~30 ;
wire \Add2~31 ;
wire \Add2~33_sumout ;
wire \Add2~34 ;
wire \Add2~35 ;
wire \Add2~37_sumout ;
wire \Add2~38 ;
wire \Add2~39 ;
wire \Add2~41_sumout ;
wire \Add2~42 ;
wire \Add2~43 ;
wire \Add2~45_sumout ;
wire \Add2~46 ;
wire \Add2~47 ;
wire \Add2~49_sumout ;
wire \Add2~50 ;
wire \Add2~51 ;
wire \Add2~53_sumout ;
wire \Add2~54 ;
wire \Add2~55 ;
wire \Add2~57_sumout ;
wire \Add2~58 ;
wire \Add2~59 ;
wire \Add2~61_sumout ;
wire \Add2~62 ;
wire \Add2~63 ;
wire \Add2~65_sumout ;
wire \Add2~66 ;
wire \Add2~67 ;
wire \Add2~69_sumout ;
wire \Add2~70 ;
wire \Add2~71 ;
wire \Add2~73_sumout ;
wire \Add2~74 ;
wire \Add2~75 ;
wire \Add2~77_sumout ;
wire \Add2~78 ;
wire \Add2~79 ;
wire \Add2~81_sumout ;
wire \Add2~82 ;
wire \Add2~83 ;
wire \Add2~85_sumout ;
wire \Add2~86 ;
wire \Add2~87 ;
wire \Add2~89_sumout ;
wire \Add2~90 ;
wire \Add2~91 ;
wire \Add2~93_sumout ;
wire \Add2~94 ;
wire \Add2~95 ;
wire \Add2~97_sumout ;
wire \Add2~98 ;
wire \Add2~99 ;
wire \Add2~101_sumout ;
wire \Add2~102 ;
wire \Add2~103 ;
wire \Add2~105_sumout ;
wire \Add2~106 ;
wire \Add2~107 ;
wire \Add2~109_sumout ;
wire \Add2~110 ;
wire \Add2~111 ;
wire \Add2~113_sumout ;
wire \Add2~114 ;
wire \Add2~115 ;
wire \Add2~117_sumout ;
wire \Add2~118 ;
wire \Add2~119 ;
wire \Add2~121_sumout ;
wire \Add2~122 ;
wire \Add2~123 ;
wire \Add2~125_sumout ;
wire \Add2~126 ;
wire \Add2~127 ;
wire \length[29]~q ;
wire \length[30]~q ;
wire \length[31]~q ;
wire \length[19]~q ;
wire \length[24]~q ;
wire \length[26]~q ;
wire \length[27]~q ;
wire \length[28]~q ;
wire \length[9]~q ;
wire \length[14]~q ;
wire \length[16]~q ;
wire \length[17]~q ;
wire \length[18]~q ;
wire \length[5]~q ;
wire \length[6]~q ;
wire \length[7]~q ;
wire \length[8]~q ;
wire \length[20]~q ;
wire \length[21]~q ;
wire \length[22]~q ;
wire \length[23]~q ;
wire \length[25]~q ;
wire \length[10]~q ;
wire \length[11]~q ;
wire \length[12]~q ;
wire \length[13]~q ;
wire \length[15]~q ;
wire \length[0]~q ;
wire \length[1]~q ;
wire \length[2]~q ;
wire \length[3]~q ;
wire \length[4]~q ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[0]~4_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[1]~8_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[2]~12_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[3]~16_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[4]~20_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[5]~24_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[6]~28_combout ;
wire \the_Computer_System_dma_2_read_data_mux|fifo_wr_data[7]~32_combout ;
wire \the_Computer_System_dma_2_read_data_mux|length_write~combout ;
wire \p1_writelength_eq_0~6_combout ;
wire \p1_writelength_eq_0~7_combout ;
wire \p1_writelength_eq_0~8_combout ;
wire \p1_done_write~1_combout ;
wire \length_eq_0~q ;
wire \p1_length_eq_0~0_combout ;
wire \p1_length_eq_0~1_combout ;
wire \p1_length_eq_0~2_combout ;
wire \p1_length_eq_0~3_combout ;
wire \p1_length_eq_0~4_combout ;
wire \p1_length_eq_0~5_combout ;
wire \p1_length_eq_0~6_combout ;
wire \p1_done_read~0_combout ;
wire \the_Computer_System_dma_2_fifo_module|p1_fifo_full~3_combout ;
wire \p1_length_eq_0~7_combout ;
wire \p1_length_eq_0~8_combout ;
wire \p1_length_eq_0~9_combout ;
wire \length_eq_0~0_combout ;
wire \length[5]~0_combout ;
wire \p1_control~0_combout ;
wire \control[12]~q ;
wire \set_software_reset_bit~0_combout ;
wire \d1_softwarereset~0_combout ;
wire \d1_softwarereset~q ;
wire \software_reset_request~0_combout ;
wire \software_reset_request~q ;
wire \reset_n~0_combout ;
wire \reset_n~q ;
wire \control[9]~q ;
wire \Add1~126 ;
wire \Add1~122 ;
wire \Add1~1_sumout ;
wire \Equal3~0_combout ;
wire \p1_writeaddress~0_combout ;
wire \writeaddress[9]~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \Add1~30 ;
wire \Add1~33_sumout ;
wire \Add1~34 ;
wire \Add1~37_sumout ;
wire \Add1~38 ;
wire \Add1~41_sumout ;
wire \Add1~42 ;
wire \Add1~45_sumout ;
wire \Add1~46 ;
wire \Add1~49_sumout ;
wire \Add1~50 ;
wire \Add1~53_sumout ;
wire \Add1~54 ;
wire \Add1~57_sumout ;
wire \Add1~58 ;
wire \Add1~61_sumout ;
wire \Add1~62 ;
wire \Add1~65_sumout ;
wire \Add1~66 ;
wire \Add1~69_sumout ;
wire \Add1~70 ;
wire \Add1~73_sumout ;
wire \Add1~74 ;
wire \Add1~77_sumout ;
wire \Add1~78 ;
wire \Add1~81_sumout ;
wire \Add1~82 ;
wire \Add1~85_sumout ;
wire \Add1~86 ;
wire \Add1~89_sumout ;
wire \Add1~90 ;
wire \Add1~93_sumout ;
wire \Add1~94 ;
wire \Add1~97_sumout ;
wire \Add1~98 ;
wire \Add1~101_sumout ;
wire \Add1~102 ;
wire \Add1~105_sumout ;
wire \Add1~106 ;
wire \Add1~109_sumout ;
wire \Add1~110 ;
wire \Add1~113_sumout ;
wire \Add1~114 ;
wire \Add1~117_sumout ;
wire \Add1~121_sumout ;
wire \Add1~125_sumout ;
wire \control[8]~q ;
wire \Add0~61_sumout ;
wire \Equal3~1_combout ;
wire \p1_readaddress~0_combout ;
wire \readaddress[13]~0_combout ;
wire \readaddress[0]~q ;
wire \Add0~62 ;
wire \Add0~57_sumout ;
wire \readaddress[1]~q ;
wire \Add0~58 ;
wire \Add0~6 ;
wire \Add0~10 ;
wire \Add0~14 ;
wire \Add0~18 ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~30 ;
wire \Add0~34 ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~46 ;
wire \Add0~50 ;
wire \Add0~54 ;
wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~9_sumout ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \Add0~29_sumout ;
wire \Add0~33_sumout ;
wire \Add0~37_sumout ;
wire \Add0~41_sumout ;
wire \Add0~45_sumout ;
wire \Add0~49_sumout ;
wire \Add0~53_sumout ;
wire \control[2]~0_combout ;
wire \Add3~113_sumout ;
wire \writelength[30]~q ;
wire \Add3~114 ;
wire \Add3~115 ;
wire \Add3~117_sumout ;
wire \writelength[1]~q ;
wire \Add3~118 ;
wire \Add3~119 ;
wire \Add3~121_sumout ;
wire \writelength[2]~q ;
wire \Add3~122 ;
wire \Add3~123 ;
wire \Add3~125_sumout ;
wire \writelength[3]~q ;
wire \Add3~126 ;
wire \Add3~127 ;
wire \Add3~49_sumout ;
wire \writelength[4]~q ;
wire \Add3~50 ;
wire \Add3~51 ;
wire \Add3~53_sumout ;
wire \writelength[5]~q ;
wire \Add3~54 ;
wire \Add3~55 ;
wire \Add3~57_sumout ;
wire \writelength[6]~q ;
wire \Add3~58 ;
wire \Add3~59 ;
wire \Add3~61_sumout ;
wire \writelength[7]~q ;
wire \Add3~62 ;
wire \Add3~63 ;
wire \Add3~65_sumout ;
wire \writelength[8]~q ;
wire \Add3~66 ;
wire \Add3~67 ;
wire \Add3~69_sumout ;
wire \writelength[9]~q ;
wire \Add3~70 ;
wire \Add3~71 ;
wire \Add3~93_sumout ;
wire \writelength[10]~q ;
wire \Add3~94 ;
wire \Add3~95 ;
wire \Add3~97_sumout ;
wire \writelength[11]~q ;
wire \Add3~98 ;
wire \Add3~99 ;
wire \Add3~101_sumout ;
wire \writelength[12]~q ;
wire \Add3~102 ;
wire \Add3~103 ;
wire \Add3~105_sumout ;
wire \writelength[13]~q ;
wire \Add3~106 ;
wire \Add3~107 ;
wire \Add3~109_sumout ;
wire \writelength[14]~q ;
wire \Add3~110 ;
wire \Add3~111 ;
wire \Add3~29_sumout ;
wire \writelength[15]~q ;
wire \Add3~30 ;
wire \Add3~31 ;
wire \Add3~33_sumout ;
wire \writelength[16]~q ;
wire \Add3~34 ;
wire \Add3~35 ;
wire \Add3~37_sumout ;
wire \writelength[17]~q ;
wire \Add3~38 ;
wire \Add3~39 ;
wire \Add3~41_sumout ;
wire \writelength[18]~q ;
wire \Add3~42 ;
wire \Add3~43 ;
wire \Add3~45_sumout ;
wire \writelength[19]~q ;
wire \Add3~46 ;
wire \Add3~47 ;
wire \Add3~73_sumout ;
wire \writelength[20]~q ;
wire \Add3~74 ;
wire \Add3~75 ;
wire \Add3~77_sumout ;
wire \writelength[21]~q ;
wire \Add3~78 ;
wire \Add3~79 ;
wire \Add3~81_sumout ;
wire \writelength[22]~q ;
wire \Add3~82 ;
wire \Add3~83 ;
wire \Add3~85_sumout ;
wire \writelength[23]~q ;
wire \Add3~86 ;
wire \Add3~87 ;
wire \Add3~89_sumout ;
wire \writelength[24]~q ;
wire \Add3~90 ;
wire \Add3~91 ;
wire \Add3~9_sumout ;
wire \writelength[25]~q ;
wire \Add3~10 ;
wire \Add3~11 ;
wire \Add3~13_sumout ;
wire \writelength[26]~q ;
wire \Add3~14 ;
wire \Add3~15 ;
wire \Add3~17_sumout ;
wire \writelength[27]~q ;
wire \Add3~18 ;
wire \Add3~19 ;
wire \Add3~21_sumout ;
wire \writelength[28]~q ;
wire \Add3~22 ;
wire \Add3~23 ;
wire \Add3~25_sumout ;
wire \writelength[29]~q ;
wire \Add3~26 ;
wire \Add3~27 ;
wire \Add3~1_sumout ;
wire \writelength[31]~q ;
wire \Add3~2 ;
wire \Add3~3 ;
wire \Add3~5_sumout ;
wire \p1_writelength_eq_0~0_combout ;
wire \p1_writelength_eq_0~1_combout ;
wire \p1_writelength_eq_0~2_combout ;
wire \p1_writelength_eq_0~3_combout ;
wire \p1_writelength_eq_0~4_combout ;
wire \p1_writelength_eq_0~5_combout ;
wire \writelength_eq_0~0_combout ;
wire \writelength_eq_0~q ;
wire \writelength[8]~0_combout ;
wire \writelength[0]~q ;
wire \Equal3~2_combout ;
wire \p1_dma_ctl_readdata[0]~0_combout ;
wire \Equal3~3_combout ;
wire \control[3]~q ;
wire \control[7]~1_combout ;
wire \control[7]~q ;
wire \p1_done_write~0_combout ;
wire \done_write~q ;
wire \done_transaction~combout ;
wire \d1_done_transaction~q ;
wire \flush_fifo~combout ;
wire \p1_readaddress~1_combout ;
wire \p1_dma_ctl_readdata~1_combout ;
wire \done~0_combout ;
wire \done~q ;
wire \p1_dma_ctl_readdata[0]~2_combout ;
wire \p1_dma_ctl_readdata[0]~combout ;
wire \p1_dma_ctl_readdata[1]~3_combout ;
wire \control[1]~q ;
wire \p1_dma_ctl_readdata[1]~4_combout ;
wire \p1_dma_ctl_readdata[1]~combout ;
wire \p1_dma_ctl_readdata[2]~43_combout ;
wire \p1_dma_ctl_readdata[3]~39_combout ;
wire \p1_dma_ctl_readdata[4]~5_combout ;
wire \control[4]~q ;
wire \len~0_combout ;
wire \len~q ;
wire \p1_dma_ctl_readdata[4]~6_combout ;
wire \p1_dma_ctl_readdata[4]~combout ;
wire \control[5]~q ;
wire \p1_dma_ctl_readdata[5]~35_combout ;
wire \control[6]~q ;
wire \p1_dma_ctl_readdata[6]~31_combout ;
wire \p1_dma_ctl_readdata[7]~27_combout ;
wire \p1_dma_ctl_readdata[8]~23_combout ;
wire \p1_dma_ctl_readdata[9]~19_combout ;
wire \control[10]~q ;
wire \p1_dma_ctl_readdata[10]~15_combout ;
wire \control[11]~q ;
wire \p1_dma_ctl_readdata[11]~11_combout ;
wire \p1_dma_ctl_readdata[12]~7_combout ;
wire \p1_dma_ctl_readdata[13]~combout ;
wire \p1_dma_ctl_readdata[14]~combout ;
wire \p1_dma_ctl_readdata[15]~combout ;
wire \Add0~2 ;
wire \Add0~65_sumout ;
wire \readaddress[16]~q ;
wire \p1_dma_ctl_readdata[16]~combout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \readaddress[17]~q ;
wire \p1_dma_ctl_readdata[17]~combout ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \readaddress[18]~q ;
wire \p1_dma_ctl_readdata[18]~combout ;
wire \Add0~74 ;
wire \Add0~77_sumout ;
wire \readaddress[19]~q ;
wire \p1_dma_ctl_readdata[19]~combout ;
wire \Add0~78 ;
wire \Add0~81_sumout ;
wire \readaddress[20]~q ;
wire \p1_dma_ctl_readdata[20]~combout ;
wire \Add0~82 ;
wire \Add0~85_sumout ;
wire \readaddress[21]~q ;
wire \p1_dma_ctl_readdata[21]~combout ;
wire \Add0~86 ;
wire \Add0~89_sumout ;
wire \readaddress[22]~q ;
wire \p1_dma_ctl_readdata[22]~combout ;
wire \Add0~90 ;
wire \Add0~93_sumout ;
wire \readaddress[23]~q ;
wire \p1_dma_ctl_readdata[23]~combout ;
wire \Add0~94 ;
wire \Add0~97_sumout ;
wire \readaddress[24]~q ;
wire \p1_dma_ctl_readdata[24]~combout ;
wire \Add0~98 ;
wire \Add0~101_sumout ;
wire \readaddress[25]~q ;
wire \p1_dma_ctl_readdata[25]~combout ;
wire \Add0~102 ;
wire \Add0~105_sumout ;
wire \readaddress[26]~q ;
wire \p1_dma_ctl_readdata[26]~combout ;
wire \Add0~106 ;
wire \Add0~109_sumout ;
wire \readaddress[27]~q ;
wire \p1_dma_ctl_readdata[27]~combout ;
wire \p1_dma_ctl_readdata[28]~combout ;
wire \p1_dma_ctl_readdata[29]~combout ;
wire \p1_dma_ctl_readdata[30]~combout ;
wire \p1_dma_ctl_readdata[31]~combout ;


Computer_System_Computer_System_dma_2_mem_write the_Computer_System_dma_2_mem_write(
	.f2h_AWREADY_0(f2h_AWREADY_0),
	.f2h_WREADY_0(f2h_WREADY_0),
	.address_taken(address_taken),
	.mem_used_7(mem_used_7),
	.src_valid(src_valid),
	.data_taken(data_taken),
	.fifo_read(fifo_read));

Computer_System_Computer_System_dma_2_mem_read the_Computer_System_dma_2_mem_read(
	.clk(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.saved_grant_0(saved_grant_0),
	.mem_used_1(mem_used_1),
	.control_3(\control[3]~q ),
	.reset_n(\reset_n~q ),
	.read_select1(read_select),
	.read_latency_shift_reg(read_latency_shift_reg),
	.control_7(\control[7]~q ),
	.p1_done_write(\p1_done_write~1_combout ),
	.p1_done_read(\p1_done_read~0_combout ),
	.p1_fifo_full(\the_Computer_System_dma_2_fifo_module|p1_fifo_full~3_combout ));

Computer_System_Computer_System_dma_2_fifo_module the_Computer_System_dma_2_fifo_module(
	.outclk_wire_0(outclk_wire_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.fifo_empty1(fifo_empty),
	.src_valid(src_valid),
	.last_write_collision1(last_write_collision),
	.last_write_data_0(last_write_data_0),
	.last_write_data_1(last_write_data_1),
	.last_write_data_2(last_write_data_2),
	.last_write_data_3(last_write_data_3),
	.last_write_data_4(last_write_data_4),
	.last_write_data_5(last_write_data_5),
	.last_write_data_6(last_write_data_6),
	.last_write_data_7(last_write_data_7),
	.last_write_data_8(last_write_data_8),
	.last_write_data_9(last_write_data_9),
	.last_write_data_10(last_write_data_10),
	.last_write_data_11(last_write_data_11),
	.last_write_data_12(last_write_data_12),
	.last_write_data_13(last_write_data_13),
	.last_write_data_14(last_write_data_14),
	.last_write_data_15(last_write_data_15),
	.last_write_data_16(last_write_data_16),
	.last_write_data_17(last_write_data_17),
	.last_write_data_18(last_write_data_18),
	.last_write_data_19(last_write_data_19),
	.last_write_data_20(last_write_data_20),
	.last_write_data_21(last_write_data_21),
	.last_write_data_22(last_write_data_22),
	.last_write_data_23(last_write_data_23),
	.last_write_data_24(last_write_data_24),
	.last_write_data_25(last_write_data_25),
	.last_write_data_26(last_write_data_26),
	.last_write_data_27(last_write_data_27),
	.last_write_data_28(last_write_data_28),
	.last_write_data_29(last_write_data_29),
	.last_write_data_30(last_write_data_30),
	.last_write_data_31(last_write_data_31),
	.fifo_read(fifo_read),
	.write_cp_ready(write_cp_ready),
	.flush_fifo(\flush_fifo~combout ),
	.src0_valid(src0_valid),
	.reset_n(\reset_n~q ),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout),
	.fifo_wr_data_0(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[0]~4_combout ),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout),
	.fifo_wr_data_1(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[1]~8_combout ),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout),
	.fifo_wr_data_2(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[2]~12_combout ),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout),
	.fifo_wr_data_3(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[3]~16_combout ),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout),
	.fifo_wr_data_4(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[4]~20_combout ),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout),
	.fifo_wr_data_5(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[5]~24_combout ),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout),
	.fifo_wr_data_6(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[6]~28_combout ),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout),
	.fifo_wr_data_7(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[7]~32_combout ),
	.l1_w8_n0_mux_dataout(l1_w8_n0_mux_dataout),
	.l1_w9_n0_mux_dataout(l1_w9_n0_mux_dataout),
	.l1_w10_n0_mux_dataout(l1_w10_n0_mux_dataout),
	.l1_w11_n0_mux_dataout(l1_w11_n0_mux_dataout),
	.l1_w12_n0_mux_dataout(l1_w12_n0_mux_dataout),
	.l1_w13_n0_mux_dataout(l1_w13_n0_mux_dataout),
	.l1_w14_n0_mux_dataout(l1_w14_n0_mux_dataout),
	.l1_w15_n0_mux_dataout(l1_w15_n0_mux_dataout),
	.l1_w24_n0_mux_dataout(l1_w24_n0_mux_dataout),
	.l1_w25_n0_mux_dataout(l1_w25_n0_mux_dataout),
	.l1_w26_n0_mux_dataout(l1_w26_n0_mux_dataout),
	.l1_w27_n0_mux_dataout(l1_w27_n0_mux_dataout),
	.l1_w28_n0_mux_dataout(l1_w28_n0_mux_dataout),
	.l1_w29_n0_mux_dataout(l1_w29_n0_mux_dataout),
	.l1_w30_n0_mux_dataout(l1_w30_n0_mux_dataout),
	.l1_w31_n0_mux_dataout(l1_w31_n0_mux_dataout),
	.read_latency_shift_reg(read_latency_shift_reg),
	.p1_fifo_full(\the_Computer_System_dma_2_fifo_module|p1_fifo_full~3_combout ));

Computer_System_Computer_System_dma_2_read_data_mux the_Computer_System_dma_2_read_data_mux(
	.ram_block1a32(ram_block1a32),
	.ram_block1a0(ram_block1a0),
	.ram_block1a33(ram_block1a33),
	.ram_block1a1(ram_block1a1),
	.ram_block1a34(ram_block1a34),
	.ram_block1a2(ram_block1a2),
	.ram_block1a35(ram_block1a35),
	.ram_block1a3(ram_block1a3),
	.ram_block1a36(ram_block1a36),
	.ram_block1a4(ram_block1a4),
	.ram_block1a37(ram_block1a37),
	.ram_block1a5(ram_block1a5),
	.ram_block1a38(ram_block1a38),
	.ram_block1a6(ram_block1a6),
	.ram_block1a39(ram_block1a39),
	.ram_block1a7(ram_block1a7),
	.ram_block1a40(ram_block1a40),
	.ram_block1a8(ram_block1a8),
	.ram_block1a41(ram_block1a41),
	.ram_block1a9(ram_block1a9),
	.ram_block1a42(ram_block1a42),
	.ram_block1a10(ram_block1a10),
	.ram_block1a43(ram_block1a43),
	.ram_block1a11(ram_block1a11),
	.ram_block1a44(ram_block1a44),
	.ram_block1a12(ram_block1a12),
	.ram_block1a45(ram_block1a45),
	.ram_block1a13(ram_block1a13),
	.ram_block1a46(ram_block1a46),
	.ram_block1a14(ram_block1a14),
	.ram_block1a47(ram_block1a47),
	.ram_block1a15(ram_block1a15),
	.ram_block1a56(ram_block1a56),
	.ram_block1a24(ram_block1a24),
	.ram_block1a57(ram_block1a57),
	.ram_block1a25(ram_block1a25),
	.ram_block1a58(ram_block1a58),
	.ram_block1a26(ram_block1a26),
	.ram_block1a59(ram_block1a59),
	.ram_block1a27(ram_block1a27),
	.ram_block1a60(ram_block1a60),
	.ram_block1a28(ram_block1a28),
	.ram_block1a61(ram_block1a61),
	.ram_block1a29(ram_block1a29),
	.ram_block1a62(ram_block1a62),
	.ram_block1a30(ram_block1a30),
	.ram_block1a63(ram_block1a63),
	.ram_block1a31(ram_block1a31),
	.clk(outclk_wire_0),
	.readaddress_0(\readaddress[0]~q ),
	.readaddress_1(\readaddress[1]~q ),
	.control_2(control_2),
	.control_0(control_0),
	.WideOr0(WideOr0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.src0_valid(src0_valid),
	.reset_n(\reset_n~q ),
	.in_data_reg_59(in_data_reg_59),
	.mem(mem),
	.in_data_reg_3(in_data_reg_3),
	.address_reg_a_0(address_reg_a_0),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout),
	.fifo_wr_data_0(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[0]~4_combout ),
	.p1_control(\p1_control~0_combout ),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout),
	.fifo_wr_data_1(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[1]~8_combout ),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout),
	.fifo_wr_data_2(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[2]~12_combout ),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout),
	.fifo_wr_data_3(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[3]~16_combout ),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout),
	.fifo_wr_data_4(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[4]~20_combout ),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout),
	.fifo_wr_data_5(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[5]~24_combout ),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout),
	.fifo_wr_data_6(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[6]~28_combout ),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout),
	.fifo_wr_data_7(\the_Computer_System_dma_2_read_data_mux|fifo_wr_data[7]~32_combout ),
	.Equal3(\Equal3~2_combout ),
	.length_write1(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.control_8(\control[8]~q ));

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(\Add2~31 ),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout(\Add2~3 ));
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~1 .shared_arith = "on";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(\Add2~3 ),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout(\Add2~7 ));
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~5 .shared_arith = "on";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(\Add2~7 ),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h000000000000FF00;
defparam \Add2~9 .shared_arith = "on";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~50 ),
	.sharein(\Add2~51 ),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout(\Add2~15 ));
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~13 .shared_arith = "on";

cyclonev_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~82 ),
	.sharein(\Add2~83 ),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout(\Add2~19 ));
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~17 .shared_arith = "on";

cyclonev_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~86 ),
	.sharein(\Add2~87 ),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout(\Add2~23 ));
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~21 .shared_arith = "on";

cyclonev_lcell_comb \Add2~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(\Add2~23 ),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(\Add2~26 ),
	.shareout(\Add2~27 ));
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~25 .shared_arith = "on";

cyclonev_lcell_comb \Add2~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~26 ),
	.sharein(\Add2~27 ),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout(\Add2~31 ));
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~29 .shared_arith = "on";

cyclonev_lcell_comb \Add2~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~66 ),
	.sharein(\Add2~67 ),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout(\Add2~35 ));
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~33 .shared_arith = "on";

cyclonev_lcell_comb \Add2~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~102 ),
	.sharein(\Add2~103 ),
	.combout(),
	.sumout(\Add2~37_sumout ),
	.cout(\Add2~38 ),
	.shareout(\Add2~39 ));
defparam \Add2~37 .extended_lut = "off";
defparam \Add2~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~37 .shared_arith = "on";

cyclonev_lcell_comb \Add2~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~106 ),
	.sharein(\Add2~107 ),
	.combout(),
	.sumout(\Add2~41_sumout ),
	.cout(\Add2~42 ),
	.shareout(\Add2~43 ));
defparam \Add2~41 .extended_lut = "off";
defparam \Add2~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~41 .shared_arith = "on";

cyclonev_lcell_comb \Add2~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~42 ),
	.sharein(\Add2~43 ),
	.combout(),
	.sumout(\Add2~45_sumout ),
	.cout(\Add2~46 ),
	.shareout(\Add2~47 ));
defparam \Add2~45 .extended_lut = "off";
defparam \Add2~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~45 .shared_arith = "on";

cyclonev_lcell_comb \Add2~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~46 ),
	.sharein(\Add2~47 ),
	.combout(),
	.sumout(\Add2~49_sumout ),
	.cout(\Add2~50 ),
	.shareout(\Add2~51 ));
defparam \Add2~49 .extended_lut = "off";
defparam \Add2~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~49 .shared_arith = "on";

cyclonev_lcell_comb \Add2~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~126 ),
	.sharein(\Add2~127 ),
	.combout(),
	.sumout(\Add2~53_sumout ),
	.cout(\Add2~54 ),
	.shareout(\Add2~55 ));
defparam \Add2~53 .extended_lut = "off";
defparam \Add2~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~53 .shared_arith = "on";

cyclonev_lcell_comb \Add2~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~54 ),
	.sharein(\Add2~55 ),
	.combout(),
	.sumout(\Add2~57_sumout ),
	.cout(\Add2~58 ),
	.shareout(\Add2~59 ));
defparam \Add2~57 .extended_lut = "off";
defparam \Add2~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~57 .shared_arith = "on";

cyclonev_lcell_comb \Add2~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~58 ),
	.sharein(\Add2~59 ),
	.combout(),
	.sumout(\Add2~61_sumout ),
	.cout(\Add2~62 ),
	.shareout(\Add2~63 ));
defparam \Add2~61 .extended_lut = "off";
defparam \Add2~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~61 .shared_arith = "on";

cyclonev_lcell_comb \Add2~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~62 ),
	.sharein(\Add2~63 ),
	.combout(),
	.sumout(\Add2~65_sumout ),
	.cout(\Add2~66 ),
	.shareout(\Add2~67 ));
defparam \Add2~65 .extended_lut = "off";
defparam \Add2~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~65 .shared_arith = "on";

cyclonev_lcell_comb \Add2~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(\Add2~15 ),
	.combout(),
	.sumout(\Add2~69_sumout ),
	.cout(\Add2~70 ),
	.shareout(\Add2~71 ));
defparam \Add2~69 .extended_lut = "off";
defparam \Add2~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~69 .shared_arith = "on";

cyclonev_lcell_comb \Add2~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~70 ),
	.sharein(\Add2~71 ),
	.combout(),
	.sumout(\Add2~73_sumout ),
	.cout(\Add2~74 ),
	.shareout(\Add2~75 ));
defparam \Add2~73 .extended_lut = "off";
defparam \Add2~73 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~73 .shared_arith = "on";

cyclonev_lcell_comb \Add2~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~74 ),
	.sharein(\Add2~75 ),
	.combout(),
	.sumout(\Add2~77_sumout ),
	.cout(\Add2~78 ),
	.shareout(\Add2~79 ));
defparam \Add2~77 .extended_lut = "off";
defparam \Add2~77 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~77 .shared_arith = "on";

cyclonev_lcell_comb \Add2~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~78 ),
	.sharein(\Add2~79 ),
	.combout(),
	.sumout(\Add2~81_sumout ),
	.cout(\Add2~82 ),
	.shareout(\Add2~83 ));
defparam \Add2~81 .extended_lut = "off";
defparam \Add2~81 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~81 .shared_arith = "on";

cyclonev_lcell_comb \Add2~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(\Add2~19 ),
	.combout(),
	.sumout(\Add2~85_sumout ),
	.cout(\Add2~86 ),
	.shareout(\Add2~87 ));
defparam \Add2~85 .extended_lut = "off";
defparam \Add2~85 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~85 .shared_arith = "on";

cyclonev_lcell_comb \Add2~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(\Add2~35 ),
	.combout(),
	.sumout(\Add2~89_sumout ),
	.cout(\Add2~90 ),
	.shareout(\Add2~91 ));
defparam \Add2~89 .extended_lut = "off";
defparam \Add2~89 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~89 .shared_arith = "on";

cyclonev_lcell_comb \Add2~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~90 ),
	.sharein(\Add2~91 ),
	.combout(),
	.sumout(\Add2~93_sumout ),
	.cout(\Add2~94 ),
	.shareout(\Add2~95 ));
defparam \Add2~93 .extended_lut = "off";
defparam \Add2~93 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~93 .shared_arith = "on";

cyclonev_lcell_comb \Add2~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~94 ),
	.sharein(\Add2~95 ),
	.combout(),
	.sumout(\Add2~97_sumout ),
	.cout(\Add2~98 ),
	.shareout(\Add2~99 ));
defparam \Add2~97 .extended_lut = "off";
defparam \Add2~97 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~97 .shared_arith = "on";

cyclonev_lcell_comb \Add2~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~98 ),
	.sharein(\Add2~99 ),
	.combout(),
	.sumout(\Add2~101_sumout ),
	.cout(\Add2~102 ),
	.shareout(\Add2~103 ));
defparam \Add2~101 .extended_lut = "off";
defparam \Add2~101 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~101 .shared_arith = "on";

cyclonev_lcell_comb \Add2~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~38 ),
	.sharein(\Add2~39 ),
	.combout(),
	.sumout(\Add2~105_sumout ),
	.cout(\Add2~106 ),
	.shareout(\Add2~107 ));
defparam \Add2~105 .extended_lut = "off";
defparam \Add2~105 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~105 .shared_arith = "on";

cyclonev_lcell_comb \Add2~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_0),
	.datad(!\length[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~109_sumout ),
	.cout(\Add2~110 ),
	.shareout(\Add2~111 ));
defparam \Add2~109 .extended_lut = "off";
defparam \Add2~109 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~109 .shared_arith = "on";

cyclonev_lcell_comb \Add2~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~110 ),
	.sharein(\Add2~111 ),
	.combout(),
	.sumout(\Add2~113_sumout ),
	.cout(\Add2~114 ),
	.shareout(\Add2~115 ));
defparam \Add2~113 .extended_lut = "off";
defparam \Add2~113 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~113 .shared_arith = "on";

cyclonev_lcell_comb \Add2~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_2),
	.datad(!\length[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~114 ),
	.sharein(\Add2~115 ),
	.combout(),
	.sumout(\Add2~117_sumout ),
	.cout(\Add2~118 ),
	.shareout(\Add2~119 ));
defparam \Add2~117 .extended_lut = "off";
defparam \Add2~117 .lut_mask = 64'h0000000F00000FF0;
defparam \Add2~117 .shared_arith = "on";

cyclonev_lcell_comb \Add2~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~118 ),
	.sharein(\Add2~119 ),
	.combout(),
	.sumout(\Add2~121_sumout ),
	.cout(\Add2~122 ),
	.shareout(\Add2~123 ));
defparam \Add2~121 .extended_lut = "off";
defparam \Add2~121 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~121 .shared_arith = "on";

cyclonev_lcell_comb \Add2~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\length[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~122 ),
	.sharein(\Add2~123 ),
	.combout(),
	.sumout(\Add2~125_sumout ),
	.cout(\Add2~126 ),
	.shareout(\Add2~127 ));
defparam \Add2~125 .extended_lut = "off";
defparam \Add2~125 .lut_mask = 64'h000000FF0000FF00;
defparam \Add2~125 .shared_arith = "on";

dffeas \length[29] (
	.clk(outclk_wire_0),
	.d(in_data_reg_29),
	.asdata(\Add2~1_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[29]~q ),
	.prn(vcc));
defparam \length[29] .is_wysiwyg = "true";
defparam \length[29] .power_up = "low";

dffeas \length[30] (
	.clk(outclk_wire_0),
	.d(in_data_reg_30),
	.asdata(\Add2~5_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[30]~q ),
	.prn(vcc));
defparam \length[30] .is_wysiwyg = "true";
defparam \length[30] .power_up = "low";

dffeas \length[31] (
	.clk(outclk_wire_0),
	.d(in_data_reg_31),
	.asdata(\Add2~9_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[31]~q ),
	.prn(vcc));
defparam \length[31] .is_wysiwyg = "true";
defparam \length[31] .power_up = "low";

dffeas \length[19] (
	.clk(outclk_wire_0),
	.d(in_data_reg_19),
	.asdata(\Add2~13_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[19]~q ),
	.prn(vcc));
defparam \length[19] .is_wysiwyg = "true";
defparam \length[19] .power_up = "low";

dffeas \length[24] (
	.clk(outclk_wire_0),
	.d(in_data_reg_24),
	.asdata(\Add2~17_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[24]~q ),
	.prn(vcc));
defparam \length[24] .is_wysiwyg = "true";
defparam \length[24] .power_up = "low";

dffeas \length[26] (
	.clk(outclk_wire_0),
	.d(in_data_reg_26),
	.asdata(\Add2~21_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[26]~q ),
	.prn(vcc));
defparam \length[26] .is_wysiwyg = "true";
defparam \length[26] .power_up = "low";

dffeas \length[27] (
	.clk(outclk_wire_0),
	.d(in_data_reg_27),
	.asdata(\Add2~25_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[27]~q ),
	.prn(vcc));
defparam \length[27] .is_wysiwyg = "true";
defparam \length[27] .power_up = "low";

dffeas \length[28] (
	.clk(outclk_wire_0),
	.d(in_data_reg_28),
	.asdata(\Add2~29_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[28]~q ),
	.prn(vcc));
defparam \length[28] .is_wysiwyg = "true";
defparam \length[28] .power_up = "low";

dffeas \length[9] (
	.clk(outclk_wire_0),
	.d(in_data_reg_9),
	.asdata(\Add2~33_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[9]~q ),
	.prn(vcc));
defparam \length[9] .is_wysiwyg = "true";
defparam \length[9] .power_up = "low";

dffeas \length[14] (
	.clk(outclk_wire_0),
	.d(in_data_reg_14),
	.asdata(\Add2~37_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[14]~q ),
	.prn(vcc));
defparam \length[14] .is_wysiwyg = "true";
defparam \length[14] .power_up = "low";

dffeas \length[16] (
	.clk(outclk_wire_0),
	.d(in_data_reg_16),
	.asdata(\Add2~41_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[16]~q ),
	.prn(vcc));
defparam \length[16] .is_wysiwyg = "true";
defparam \length[16] .power_up = "low";

dffeas \length[17] (
	.clk(outclk_wire_0),
	.d(in_data_reg_17),
	.asdata(\Add2~45_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[17]~q ),
	.prn(vcc));
defparam \length[17] .is_wysiwyg = "true";
defparam \length[17] .power_up = "low";

dffeas \length[18] (
	.clk(outclk_wire_0),
	.d(in_data_reg_18),
	.asdata(\Add2~49_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[18]~q ),
	.prn(vcc));
defparam \length[18] .is_wysiwyg = "true";
defparam \length[18] .power_up = "low";

dffeas \length[5] (
	.clk(outclk_wire_0),
	.d(in_data_reg_5),
	.asdata(\Add2~53_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[5]~q ),
	.prn(vcc));
defparam \length[5] .is_wysiwyg = "true";
defparam \length[5] .power_up = "low";

dffeas \length[6] (
	.clk(outclk_wire_0),
	.d(in_data_reg_6),
	.asdata(\Add2~57_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[6]~q ),
	.prn(vcc));
defparam \length[6] .is_wysiwyg = "true";
defparam \length[6] .power_up = "low";

dffeas \length[7] (
	.clk(outclk_wire_0),
	.d(in_data_reg_7),
	.asdata(\Add2~61_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[7]~q ),
	.prn(vcc));
defparam \length[7] .is_wysiwyg = "true";
defparam \length[7] .power_up = "low";

dffeas \length[8] (
	.clk(outclk_wire_0),
	.d(in_data_reg_8),
	.asdata(\Add2~65_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[8]~q ),
	.prn(vcc));
defparam \length[8] .is_wysiwyg = "true";
defparam \length[8] .power_up = "low";

dffeas \length[20] (
	.clk(outclk_wire_0),
	.d(in_data_reg_20),
	.asdata(\Add2~69_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[20]~q ),
	.prn(vcc));
defparam \length[20] .is_wysiwyg = "true";
defparam \length[20] .power_up = "low";

dffeas \length[21] (
	.clk(outclk_wire_0),
	.d(in_data_reg_21),
	.asdata(\Add2~73_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[21]~q ),
	.prn(vcc));
defparam \length[21] .is_wysiwyg = "true";
defparam \length[21] .power_up = "low";

dffeas \length[22] (
	.clk(outclk_wire_0),
	.d(in_data_reg_22),
	.asdata(\Add2~77_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[22]~q ),
	.prn(vcc));
defparam \length[22] .is_wysiwyg = "true";
defparam \length[22] .power_up = "low";

dffeas \length[23] (
	.clk(outclk_wire_0),
	.d(in_data_reg_23),
	.asdata(\Add2~81_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[23]~q ),
	.prn(vcc));
defparam \length[23] .is_wysiwyg = "true";
defparam \length[23] .power_up = "low";

dffeas \length[25] (
	.clk(outclk_wire_0),
	.d(in_data_reg_25),
	.asdata(\Add2~85_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[25]~q ),
	.prn(vcc));
defparam \length[25] .is_wysiwyg = "true";
defparam \length[25] .power_up = "low";

dffeas \length[10] (
	.clk(outclk_wire_0),
	.d(in_data_reg_10),
	.asdata(\Add2~89_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[10]~q ),
	.prn(vcc));
defparam \length[10] .is_wysiwyg = "true";
defparam \length[10] .power_up = "low";

dffeas \length[11] (
	.clk(outclk_wire_0),
	.d(in_data_reg_11),
	.asdata(\Add2~93_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[11]~q ),
	.prn(vcc));
defparam \length[11] .is_wysiwyg = "true";
defparam \length[11] .power_up = "low";

dffeas \length[12] (
	.clk(outclk_wire_0),
	.d(in_data_reg_12),
	.asdata(\Add2~97_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[12]~q ),
	.prn(vcc));
defparam \length[12] .is_wysiwyg = "true";
defparam \length[12] .power_up = "low";

dffeas \length[13] (
	.clk(outclk_wire_0),
	.d(in_data_reg_13),
	.asdata(\Add2~101_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[13]~q ),
	.prn(vcc));
defparam \length[13] .is_wysiwyg = "true";
defparam \length[13] .power_up = "low";

dffeas \length[15] (
	.clk(outclk_wire_0),
	.d(in_data_reg_15),
	.asdata(\Add2~105_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[15]~q ),
	.prn(vcc));
defparam \length[15] .is_wysiwyg = "true";
defparam \length[15] .power_up = "low";

dffeas \length[0] (
	.clk(outclk_wire_0),
	.d(in_data_reg_0),
	.asdata(\Add2~109_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[0]~q ),
	.prn(vcc));
defparam \length[0] .is_wysiwyg = "true";
defparam \length[0] .power_up = "low";

dffeas \length[1] (
	.clk(outclk_wire_0),
	.d(in_data_reg_1),
	.asdata(\Add2~113_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[1]~q ),
	.prn(vcc));
defparam \length[1] .is_wysiwyg = "true";
defparam \length[1] .power_up = "low";

dffeas \length[2] (
	.clk(outclk_wire_0),
	.d(in_data_reg_2),
	.asdata(\Add2~117_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[2]~q ),
	.prn(vcc));
defparam \length[2] .is_wysiwyg = "true";
defparam \length[2] .power_up = "low";

dffeas \length[3] (
	.clk(outclk_wire_0),
	.d(in_data_reg_3),
	.asdata(\Add2~121_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[3]~q ),
	.prn(vcc));
defparam \length[3] .is_wysiwyg = "true";
defparam \length[3] .power_up = "low";

dffeas \length[4] (
	.clk(outclk_wire_0),
	.d(in_data_reg_4),
	.asdata(\Add2~125_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\length[5]~0_combout ),
	.q(\length[4]~q ),
	.prn(vcc));
defparam \length[4] .is_wysiwyg = "true";
defparam \length[4] .power_up = "low";

cyclonev_lcell_comb \p1_writelength_eq_0~6 (
	.dataa(!\Add3~49_sumout ),
	.datab(!\Add3~53_sumout ),
	.datac(!\Add3~57_sumout ),
	.datad(!\Add3~61_sumout ),
	.datae(!\Add3~65_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~6 .extended_lut = "off";
defparam \p1_writelength_eq_0~6 .lut_mask = 64'h8000000080000000;
defparam \p1_writelength_eq_0~6 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~7 (
	.dataa(!\Add3~69_sumout ),
	.datab(!\Add3~29_sumout ),
	.datac(!\Add3~33_sumout ),
	.datad(!\Add3~37_sumout ),
	.datae(!\Add3~41_sumout ),
	.dataf(!\p1_writelength_eq_0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~7 .extended_lut = "off";
defparam \p1_writelength_eq_0~7 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~7 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~8 (
	.dataa(!\Add3~45_sumout ),
	.datab(!\Add3~9_sumout ),
	.datac(!\Add3~13_sumout ),
	.datad(!\Add3~17_sumout ),
	.datae(!\Add3~21_sumout ),
	.dataf(!\p1_writelength_eq_0~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~8 .extended_lut = "off";
defparam \p1_writelength_eq_0~8 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~8 .shared_arith = "off";

cyclonev_lcell_comb \p1_done_write~1 (
	.dataa(!\writelength_eq_0~q ),
	.datab(!\Add3~25_sumout ),
	.datac(!\Add3~1_sumout ),
	.datad(!\Add3~5_sumout ),
	.datae(!\p1_writelength_eq_0~8_combout ),
	.dataf(!\p1_writelength_eq_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_done_write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_done_write~1 .extended_lut = "off";
defparam \p1_done_write~1 .lut_mask = 64'hAAAAAAAAAAAAEAAA;
defparam \p1_done_write~1 .shared_arith = "off";

dffeas length_eq_0(
	.clk(outclk_wire_0),
	.d(\length_eq_0~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\length_eq_0~q ),
	.prn(vcc));
defparam length_eq_0.is_wysiwyg = "true";
defparam length_eq_0.power_up = "low";

cyclonev_lcell_comb \p1_length_eq_0~0 (
	.dataa(!\Add2~53_sumout ),
	.datab(!\Add2~57_sumout ),
	.datac(!\Add2~61_sumout ),
	.datad(!\Add2~65_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~0 .extended_lut = "off";
defparam \p1_length_eq_0~0 .lut_mask = 64'h8000800080008000;
defparam \p1_length_eq_0~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~1 (
	.dataa(!\Add2~33_sumout ),
	.datab(!\Add2~37_sumout ),
	.datac(!\Add2~41_sumout ),
	.datad(!\Add2~45_sumout ),
	.datae(!\Add2~49_sumout ),
	.dataf(!\p1_length_eq_0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~1 .extended_lut = "off";
defparam \p1_length_eq_0~1 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~2 (
	.dataa(!\Add2~13_sumout ),
	.datab(!\Add2~17_sumout ),
	.datac(!\Add2~21_sumout ),
	.datad(!\Add2~25_sumout ),
	.datae(!\Add2~29_sumout ),
	.dataf(!\p1_length_eq_0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~2 .extended_lut = "off";
defparam \p1_length_eq_0~2 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~3 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!read_select),
	.datae(!\length_eq_0~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~3 .extended_lut = "off";
defparam \p1_length_eq_0~3 .lut_mask = 64'h0000001000000010;
defparam \p1_length_eq_0~3 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~4 (
	.dataa(!\Add2~109_sumout ),
	.datab(!\Add2~113_sumout ),
	.datac(!\Add2~117_sumout ),
	.datad(!\Add2~121_sumout ),
	.datae(!\Add2~125_sumout ),
	.dataf(!\p1_length_eq_0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~4 .extended_lut = "off";
defparam \p1_length_eq_0~4 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~4 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~5 (
	.dataa(!\Add2~89_sumout ),
	.datab(!\Add2~93_sumout ),
	.datac(!\Add2~97_sumout ),
	.datad(!\Add2~101_sumout ),
	.datae(!\Add2~105_sumout ),
	.dataf(!\p1_length_eq_0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~5 .extended_lut = "off";
defparam \p1_length_eq_0~5 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~5 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~6 (
	.dataa(!\Add2~69_sumout ),
	.datab(!\Add2~73_sumout ),
	.datac(!\Add2~77_sumout ),
	.datad(!\Add2~81_sumout ),
	.datae(!\Add2~85_sumout ),
	.dataf(!\p1_length_eq_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~6 .extended_lut = "off";
defparam \p1_length_eq_0~6 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~6 .shared_arith = "off";

cyclonev_lcell_comb \p1_done_read~0 (
	.dataa(!\length_eq_0~q ),
	.datab(!\Add2~1_sumout ),
	.datac(!\Add2~5_sumout ),
	.datad(!\Add2~9_sumout ),
	.datae(!\p1_length_eq_0~2_combout ),
	.dataf(!\p1_length_eq_0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_done_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_done_read~0 .extended_lut = "off";
defparam \p1_done_read~0 .lut_mask = 64'h5555555555551555;
defparam \p1_done_read~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~7 (
	.dataa(!\Add2~53_sumout ),
	.datab(!\Add2~57_sumout ),
	.datac(!\Add2~61_sumout ),
	.datad(!\Add2~65_sumout ),
	.datae(!\Add2~33_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~7 .extended_lut = "off";
defparam \p1_length_eq_0~7 .lut_mask = 64'h8000000080000000;
defparam \p1_length_eq_0~7 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~8 (
	.dataa(!\Add2~37_sumout ),
	.datab(!\Add2~41_sumout ),
	.datac(!\Add2~45_sumout ),
	.datad(!\Add2~49_sumout ),
	.datae(!\Add2~13_sumout ),
	.dataf(!\p1_length_eq_0~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~8 .extended_lut = "off";
defparam \p1_length_eq_0~8 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~8 .shared_arith = "off";

cyclonev_lcell_comb \p1_length_eq_0~9 (
	.dataa(!\Add2~17_sumout ),
	.datab(!\Add2~21_sumout ),
	.datac(!\Add2~25_sumout ),
	.datad(!\Add2~29_sumout ),
	.datae(!\Add2~1_sumout ),
	.dataf(!\p1_length_eq_0~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_length_eq_0~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_length_eq_0~9 .extended_lut = "off";
defparam \p1_length_eq_0~9 .lut_mask = 64'h0000000080000000;
defparam \p1_length_eq_0~9 .shared_arith = "off";

cyclonev_lcell_comb \length_eq_0~0 (
	.dataa(!\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.datab(!\length_eq_0~q ),
	.datac(!\Add2~5_sumout ),
	.datad(!\Add2~9_sumout ),
	.datae(!\p1_length_eq_0~9_combout ),
	.dataf(!\p1_length_eq_0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\length_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \length_eq_0~0 .extended_lut = "off";
defparam \length_eq_0~0 .lut_mask = 64'hBBBBBBBBBBBBABBB;
defparam \length_eq_0~0 .shared_arith = "off";

cyclonev_lcell_comb \length[5]~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~2_combout ),
	.dataf(!\p1_length_eq_0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\length[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \length[5]~0 .extended_lut = "off";
defparam \length[5]~0 .lut_mask = 64'h00000008FFFFFFFF;
defparam \length[5]~0 .shared_arith = "off";

dffeas \writeaddress[2] (
	.clk(outclk_wire_0),
	.d(\Add1~1_sumout ),
	.asdata(in_data_reg_2),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_2),
	.prn(vcc));
defparam \writeaddress[2] .is_wysiwyg = "true";
defparam \writeaddress[2] .power_up = "low";

dffeas \writeaddress[3] (
	.clk(outclk_wire_0),
	.d(\Add1~5_sumout ),
	.asdata(in_data_reg_3),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_3),
	.prn(vcc));
defparam \writeaddress[3] .is_wysiwyg = "true";
defparam \writeaddress[3] .power_up = "low";

dffeas \writeaddress[4] (
	.clk(outclk_wire_0),
	.d(\Add1~9_sumout ),
	.asdata(in_data_reg_4),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_4),
	.prn(vcc));
defparam \writeaddress[4] .is_wysiwyg = "true";
defparam \writeaddress[4] .power_up = "low";

dffeas \writeaddress[5] (
	.clk(outclk_wire_0),
	.d(\Add1~13_sumout ),
	.asdata(in_data_reg_5),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_5),
	.prn(vcc));
defparam \writeaddress[5] .is_wysiwyg = "true";
defparam \writeaddress[5] .power_up = "low";

dffeas \writeaddress[6] (
	.clk(outclk_wire_0),
	.d(\Add1~17_sumout ),
	.asdata(in_data_reg_6),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_6),
	.prn(vcc));
defparam \writeaddress[6] .is_wysiwyg = "true";
defparam \writeaddress[6] .power_up = "low";

dffeas \writeaddress[7] (
	.clk(outclk_wire_0),
	.d(\Add1~21_sumout ),
	.asdata(in_data_reg_7),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_7),
	.prn(vcc));
defparam \writeaddress[7] .is_wysiwyg = "true";
defparam \writeaddress[7] .power_up = "low";

dffeas \writeaddress[8] (
	.clk(outclk_wire_0),
	.d(\Add1~25_sumout ),
	.asdata(in_data_reg_8),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_8),
	.prn(vcc));
defparam \writeaddress[8] .is_wysiwyg = "true";
defparam \writeaddress[8] .power_up = "low";

dffeas \writeaddress[9] (
	.clk(outclk_wire_0),
	.d(\Add1~29_sumout ),
	.asdata(in_data_reg_9),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_9),
	.prn(vcc));
defparam \writeaddress[9] .is_wysiwyg = "true";
defparam \writeaddress[9] .power_up = "low";

dffeas \writeaddress[10] (
	.clk(outclk_wire_0),
	.d(\Add1~33_sumout ),
	.asdata(in_data_reg_10),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_10),
	.prn(vcc));
defparam \writeaddress[10] .is_wysiwyg = "true";
defparam \writeaddress[10] .power_up = "low";

dffeas \writeaddress[11] (
	.clk(outclk_wire_0),
	.d(\Add1~37_sumout ),
	.asdata(in_data_reg_11),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_11),
	.prn(vcc));
defparam \writeaddress[11] .is_wysiwyg = "true";
defparam \writeaddress[11] .power_up = "low";

dffeas \writeaddress[12] (
	.clk(outclk_wire_0),
	.d(\Add1~41_sumout ),
	.asdata(in_data_reg_12),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_12),
	.prn(vcc));
defparam \writeaddress[12] .is_wysiwyg = "true";
defparam \writeaddress[12] .power_up = "low";

dffeas \writeaddress[13] (
	.clk(outclk_wire_0),
	.d(\Add1~45_sumout ),
	.asdata(in_data_reg_13),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_13),
	.prn(vcc));
defparam \writeaddress[13] .is_wysiwyg = "true";
defparam \writeaddress[13] .power_up = "low";

dffeas \writeaddress[14] (
	.clk(outclk_wire_0),
	.d(\Add1~49_sumout ),
	.asdata(in_data_reg_14),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_14),
	.prn(vcc));
defparam \writeaddress[14] .is_wysiwyg = "true";
defparam \writeaddress[14] .power_up = "low";

dffeas \writeaddress[15] (
	.clk(outclk_wire_0),
	.d(\Add1~53_sumout ),
	.asdata(in_data_reg_15),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_15),
	.prn(vcc));
defparam \writeaddress[15] .is_wysiwyg = "true";
defparam \writeaddress[15] .power_up = "low";

dffeas \writeaddress[16] (
	.clk(outclk_wire_0),
	.d(\Add1~57_sumout ),
	.asdata(in_data_reg_16),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_16),
	.prn(vcc));
defparam \writeaddress[16] .is_wysiwyg = "true";
defparam \writeaddress[16] .power_up = "low";

dffeas \writeaddress[17] (
	.clk(outclk_wire_0),
	.d(\Add1~61_sumout ),
	.asdata(in_data_reg_17),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_17),
	.prn(vcc));
defparam \writeaddress[17] .is_wysiwyg = "true";
defparam \writeaddress[17] .power_up = "low";

dffeas \writeaddress[18] (
	.clk(outclk_wire_0),
	.d(\Add1~65_sumout ),
	.asdata(in_data_reg_18),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_18),
	.prn(vcc));
defparam \writeaddress[18] .is_wysiwyg = "true";
defparam \writeaddress[18] .power_up = "low";

dffeas \writeaddress[19] (
	.clk(outclk_wire_0),
	.d(\Add1~69_sumout ),
	.asdata(in_data_reg_19),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_19),
	.prn(vcc));
defparam \writeaddress[19] .is_wysiwyg = "true";
defparam \writeaddress[19] .power_up = "low";

dffeas \writeaddress[20] (
	.clk(outclk_wire_0),
	.d(\Add1~73_sumout ),
	.asdata(in_data_reg_20),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_20),
	.prn(vcc));
defparam \writeaddress[20] .is_wysiwyg = "true";
defparam \writeaddress[20] .power_up = "low";

dffeas \writeaddress[21] (
	.clk(outclk_wire_0),
	.d(\Add1~77_sumout ),
	.asdata(in_data_reg_21),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_21),
	.prn(vcc));
defparam \writeaddress[21] .is_wysiwyg = "true";
defparam \writeaddress[21] .power_up = "low";

dffeas \writeaddress[22] (
	.clk(outclk_wire_0),
	.d(\Add1~81_sumout ),
	.asdata(in_data_reg_22),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_22),
	.prn(vcc));
defparam \writeaddress[22] .is_wysiwyg = "true";
defparam \writeaddress[22] .power_up = "low";

dffeas \writeaddress[23] (
	.clk(outclk_wire_0),
	.d(\Add1~85_sumout ),
	.asdata(in_data_reg_23),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_23),
	.prn(vcc));
defparam \writeaddress[23] .is_wysiwyg = "true";
defparam \writeaddress[23] .power_up = "low";

dffeas \writeaddress[24] (
	.clk(outclk_wire_0),
	.d(\Add1~89_sumout ),
	.asdata(in_data_reg_24),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_24),
	.prn(vcc));
defparam \writeaddress[24] .is_wysiwyg = "true";
defparam \writeaddress[24] .power_up = "low";

dffeas \writeaddress[25] (
	.clk(outclk_wire_0),
	.d(\Add1~93_sumout ),
	.asdata(in_data_reg_25),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_25),
	.prn(vcc));
defparam \writeaddress[25] .is_wysiwyg = "true";
defparam \writeaddress[25] .power_up = "low";

dffeas \writeaddress[26] (
	.clk(outclk_wire_0),
	.d(\Add1~97_sumout ),
	.asdata(in_data_reg_26),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_26),
	.prn(vcc));
defparam \writeaddress[26] .is_wysiwyg = "true";
defparam \writeaddress[26] .power_up = "low";

dffeas \writeaddress[27] (
	.clk(outclk_wire_0),
	.d(\Add1~101_sumout ),
	.asdata(in_data_reg_27),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_27),
	.prn(vcc));
defparam \writeaddress[27] .is_wysiwyg = "true";
defparam \writeaddress[27] .power_up = "low";

dffeas \writeaddress[28] (
	.clk(outclk_wire_0),
	.d(\Add1~105_sumout ),
	.asdata(in_data_reg_28),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_28),
	.prn(vcc));
defparam \writeaddress[28] .is_wysiwyg = "true";
defparam \writeaddress[28] .power_up = "low";

dffeas \writeaddress[29] (
	.clk(outclk_wire_0),
	.d(\Add1~109_sumout ),
	.asdata(in_data_reg_29),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_29),
	.prn(vcc));
defparam \writeaddress[29] .is_wysiwyg = "true";
defparam \writeaddress[29] .power_up = "low";

dffeas \writeaddress[30] (
	.clk(outclk_wire_0),
	.d(\Add1~113_sumout ),
	.asdata(in_data_reg_30),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_30),
	.prn(vcc));
defparam \writeaddress[30] .is_wysiwyg = "true";
defparam \writeaddress[30] .power_up = "low";

dffeas \writeaddress[31] (
	.clk(outclk_wire_0),
	.d(\Add1~117_sumout ),
	.asdata(in_data_reg_31),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_31),
	.prn(vcc));
defparam \writeaddress[31] .is_wysiwyg = "true";
defparam \writeaddress[31] .power_up = "low";

dffeas \writeaddress[1] (
	.clk(outclk_wire_0),
	.d(\Add1~121_sumout ),
	.asdata(in_data_reg_1),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_1),
	.prn(vcc));
defparam \writeaddress[1] .is_wysiwyg = "true";
defparam \writeaddress[1] .power_up = "low";

dffeas \writeaddress[0] (
	.clk(outclk_wire_0),
	.d(\Add1~125_sumout ),
	.asdata(in_data_reg_0),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_writeaddress~0_combout ),
	.ena(\writeaddress[9]~0_combout ),
	.q(writeaddress_0),
	.prn(vcc));
defparam \writeaddress[0] .is_wysiwyg = "true";
defparam \writeaddress[0] .power_up = "low";

dffeas \readaddress[15] (
	.clk(outclk_wire_0),
	.d(\Add0~1_sumout ),
	.asdata(in_data_reg_15),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_15),
	.prn(vcc));
defparam \readaddress[15] .is_wysiwyg = "true";
defparam \readaddress[15] .power_up = "low";

dffeas \readaddress[2] (
	.clk(outclk_wire_0),
	.d(\Add0~5_sumout ),
	.asdata(in_data_reg_2),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_2),
	.prn(vcc));
defparam \readaddress[2] .is_wysiwyg = "true";
defparam \readaddress[2] .power_up = "low";

dffeas \readaddress[3] (
	.clk(outclk_wire_0),
	.d(\Add0~9_sumout ),
	.asdata(in_data_reg_3),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_3),
	.prn(vcc));
defparam \readaddress[3] .is_wysiwyg = "true";
defparam \readaddress[3] .power_up = "low";

dffeas \readaddress[4] (
	.clk(outclk_wire_0),
	.d(\Add0~13_sumout ),
	.asdata(in_data_reg_4),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_4),
	.prn(vcc));
defparam \readaddress[4] .is_wysiwyg = "true";
defparam \readaddress[4] .power_up = "low";

dffeas \readaddress[5] (
	.clk(outclk_wire_0),
	.d(\Add0~17_sumout ),
	.asdata(in_data_reg_5),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_5),
	.prn(vcc));
defparam \readaddress[5] .is_wysiwyg = "true";
defparam \readaddress[5] .power_up = "low";

dffeas \readaddress[6] (
	.clk(outclk_wire_0),
	.d(\Add0~21_sumout ),
	.asdata(in_data_reg_6),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_6),
	.prn(vcc));
defparam \readaddress[6] .is_wysiwyg = "true";
defparam \readaddress[6] .power_up = "low";

dffeas \readaddress[7] (
	.clk(outclk_wire_0),
	.d(\Add0~25_sumout ),
	.asdata(in_data_reg_7),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_7),
	.prn(vcc));
defparam \readaddress[7] .is_wysiwyg = "true";
defparam \readaddress[7] .power_up = "low";

dffeas \readaddress[8] (
	.clk(outclk_wire_0),
	.d(\Add0~29_sumout ),
	.asdata(in_data_reg_8),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_8),
	.prn(vcc));
defparam \readaddress[8] .is_wysiwyg = "true";
defparam \readaddress[8] .power_up = "low";

dffeas \readaddress[9] (
	.clk(outclk_wire_0),
	.d(\Add0~33_sumout ),
	.asdata(in_data_reg_9),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_9),
	.prn(vcc));
defparam \readaddress[9] .is_wysiwyg = "true";
defparam \readaddress[9] .power_up = "low";

dffeas \readaddress[10] (
	.clk(outclk_wire_0),
	.d(\Add0~37_sumout ),
	.asdata(in_data_reg_10),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_10),
	.prn(vcc));
defparam \readaddress[10] .is_wysiwyg = "true";
defparam \readaddress[10] .power_up = "low";

dffeas \readaddress[11] (
	.clk(outclk_wire_0),
	.d(\Add0~41_sumout ),
	.asdata(in_data_reg_11),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_11),
	.prn(vcc));
defparam \readaddress[11] .is_wysiwyg = "true";
defparam \readaddress[11] .power_up = "low";

dffeas \readaddress[12] (
	.clk(outclk_wire_0),
	.d(\Add0~45_sumout ),
	.asdata(in_data_reg_12),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_12),
	.prn(vcc));
defparam \readaddress[12] .is_wysiwyg = "true";
defparam \readaddress[12] .power_up = "low";

dffeas \readaddress[13] (
	.clk(outclk_wire_0),
	.d(\Add0~49_sumout ),
	.asdata(in_data_reg_13),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_13),
	.prn(vcc));
defparam \readaddress[13] .is_wysiwyg = "true";
defparam \readaddress[13] .power_up = "low";

dffeas \readaddress[14] (
	.clk(outclk_wire_0),
	.d(\Add0~53_sumout ),
	.asdata(in_data_reg_14),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(readaddress_14),
	.prn(vcc));
defparam \readaddress[14] .is_wysiwyg = "true";
defparam \readaddress[14] .power_up = "low";

dffeas \control[2] (
	.clk(outclk_wire_0),
	.d(\control[2]~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(control_2),
	.prn(vcc));
defparam \control[2] .is_wysiwyg = "true";
defparam \control[2] .power_up = "low";

dffeas \control[0] (
	.clk(outclk_wire_0),
	.d(in_data_reg_0),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(control_0),
	.prn(vcc));
defparam \control[0] .is_wysiwyg = "true";
defparam \control[0] .power_up = "low";

cyclonev_lcell_comb \write_writedata~0 (
	.dataa(!last_write_collision),
	.datab(!last_write_data_0),
	.datac(!q_b_0),
	.datad(!control_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~0 .extended_lut = "off";
defparam \write_writedata~0 .lut_mask = 64'h001B001B001B001B;
defparam \write_writedata~0 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~1 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_1),
	.datad(!q_b_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~1 .extended_lut = "off";
defparam \write_writedata~1 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~1 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~2 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_2),
	.datad(!q_b_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata2),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~2 .extended_lut = "off";
defparam \write_writedata~2 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~2 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~3 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_3),
	.datad(!q_b_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata3),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~3 .extended_lut = "off";
defparam \write_writedata~3 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~3 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~4 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_4),
	.datad(!q_b_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata4),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~4 .extended_lut = "off";
defparam \write_writedata~4 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~4 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~5 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_5),
	.datad(!q_b_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata5),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~5 .extended_lut = "off";
defparam \write_writedata~5 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~5 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~6 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_6),
	.datad(!q_b_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata6),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~6 .extended_lut = "off";
defparam \write_writedata~6 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~6 .shared_arith = "off";

cyclonev_lcell_comb \write_writedata~7 (
	.dataa(!last_write_collision),
	.datab(!control_0),
	.datac(!last_write_data_7),
	.datad(!q_b_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_writedata7),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_writedata~7 .extended_lut = "off";
defparam \write_writedata~7 .lut_mask = 64'h0123012301230123;
defparam \write_writedata~7 .shared_arith = "off";

dffeas \dma_ctl_readdata[0] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[0]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_0),
	.prn(vcc));
defparam \dma_ctl_readdata[0] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[0] .power_up = "low";

dffeas \dma_ctl_readdata[1] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[1]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_1),
	.prn(vcc));
defparam \dma_ctl_readdata[1] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[1] .power_up = "low";

dffeas \dma_ctl_readdata[2] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[2]~43_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_2),
	.prn(vcc));
defparam \dma_ctl_readdata[2] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[2] .power_up = "low";

dffeas \dma_ctl_readdata[3] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[3]~39_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_3),
	.prn(vcc));
defparam \dma_ctl_readdata[3] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[3] .power_up = "low";

dffeas \dma_ctl_readdata[4] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[4]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_4),
	.prn(vcc));
defparam \dma_ctl_readdata[4] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[4] .power_up = "low";

dffeas \dma_ctl_readdata[5] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[5]~35_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_5),
	.prn(vcc));
defparam \dma_ctl_readdata[5] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[5] .power_up = "low";

dffeas \dma_ctl_readdata[6] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[6]~31_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_6),
	.prn(vcc));
defparam \dma_ctl_readdata[6] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[6] .power_up = "low";

dffeas \dma_ctl_readdata[7] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[7]~27_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_7),
	.prn(vcc));
defparam \dma_ctl_readdata[7] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[7] .power_up = "low";

dffeas \dma_ctl_readdata[8] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[8]~23_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_8),
	.prn(vcc));
defparam \dma_ctl_readdata[8] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[8] .power_up = "low";

dffeas \dma_ctl_readdata[9] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[9]~19_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_9),
	.prn(vcc));
defparam \dma_ctl_readdata[9] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[9] .power_up = "low";

dffeas \dma_ctl_readdata[10] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[10]~15_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_10),
	.prn(vcc));
defparam \dma_ctl_readdata[10] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[10] .power_up = "low";

dffeas \dma_ctl_readdata[11] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[11]~11_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_11),
	.prn(vcc));
defparam \dma_ctl_readdata[11] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[11] .power_up = "low";

dffeas \dma_ctl_readdata[12] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[12]~7_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_12),
	.prn(vcc));
defparam \dma_ctl_readdata[12] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[12] .power_up = "low";

dffeas \dma_ctl_readdata[13] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[13]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_13),
	.prn(vcc));
defparam \dma_ctl_readdata[13] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[13] .power_up = "low";

dffeas \dma_ctl_readdata[14] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[14]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_14),
	.prn(vcc));
defparam \dma_ctl_readdata[14] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[14] .power_up = "low";

dffeas \dma_ctl_readdata[15] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[15]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_15),
	.prn(vcc));
defparam \dma_ctl_readdata[15] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[15] .power_up = "low";

dffeas \dma_ctl_readdata[16] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[16]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_16),
	.prn(vcc));
defparam \dma_ctl_readdata[16] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[16] .power_up = "low";

dffeas \dma_ctl_readdata[17] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[17]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_17),
	.prn(vcc));
defparam \dma_ctl_readdata[17] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[17] .power_up = "low";

dffeas \dma_ctl_readdata[18] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[18]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_18),
	.prn(vcc));
defparam \dma_ctl_readdata[18] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[18] .power_up = "low";

dffeas \dma_ctl_readdata[19] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[19]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_19),
	.prn(vcc));
defparam \dma_ctl_readdata[19] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[19] .power_up = "low";

dffeas \dma_ctl_readdata[20] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[20]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_20),
	.prn(vcc));
defparam \dma_ctl_readdata[20] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[20] .power_up = "low";

dffeas \dma_ctl_readdata[21] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[21]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_21),
	.prn(vcc));
defparam \dma_ctl_readdata[21] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[21] .power_up = "low";

dffeas \dma_ctl_readdata[22] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[22]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_22),
	.prn(vcc));
defparam \dma_ctl_readdata[22] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[22] .power_up = "low";

dffeas \dma_ctl_readdata[23] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[23]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_23),
	.prn(vcc));
defparam \dma_ctl_readdata[23] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[23] .power_up = "low";

dffeas \dma_ctl_readdata[24] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[24]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_24),
	.prn(vcc));
defparam \dma_ctl_readdata[24] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[24] .power_up = "low";

dffeas \dma_ctl_readdata[25] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[25]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_25),
	.prn(vcc));
defparam \dma_ctl_readdata[25] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[25] .power_up = "low";

dffeas \dma_ctl_readdata[26] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[26]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_26),
	.prn(vcc));
defparam \dma_ctl_readdata[26] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[26] .power_up = "low";

dffeas \dma_ctl_readdata[27] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[27]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_27),
	.prn(vcc));
defparam \dma_ctl_readdata[27] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[27] .power_up = "low";

dffeas \dma_ctl_readdata[28] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[28]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_28),
	.prn(vcc));
defparam \dma_ctl_readdata[28] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[28] .power_up = "low";

dffeas \dma_ctl_readdata[29] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[29]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_29),
	.prn(vcc));
defparam \dma_ctl_readdata[29] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[29] .power_up = "low";

dffeas \dma_ctl_readdata[30] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[30]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_30),
	.prn(vcc));
defparam \dma_ctl_readdata[30] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[30] .power_up = "low";

dffeas \dma_ctl_readdata[31] (
	.clk(outclk_wire_0),
	.d(\p1_dma_ctl_readdata[31]~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dma_ctl_readdata_31),
	.prn(vcc));
defparam \dma_ctl_readdata[31] .is_wysiwyg = "true";
defparam \dma_ctl_readdata[31] .power_up = "low";

cyclonev_lcell_comb \p1_control~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!int_nxt_addr_reg_dly_4),
	.dataf(!int_nxt_addr_reg_dly_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_control~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_control~0 .extended_lut = "off";
defparam \p1_control~0 .lut_mask = 64'h0000000000000008;
defparam \p1_control~0 .shared_arith = "off";

dffeas \control[12] (
	.clk(outclk_wire_0),
	.d(in_data_reg_12),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[12]~q ),
	.prn(vcc));
defparam \control[12] .is_wysiwyg = "true";
defparam \control[12] .power_up = "low";

cyclonev_lcell_comb \set_software_reset_bit~0 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!in_data_reg_12),
	.datae(!\p1_control~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\set_software_reset_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \set_software_reset_bit~0 .extended_lut = "off";
defparam \set_software_reset_bit~0 .lut_mask = 64'h000000FE000000FE;
defparam \set_software_reset_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \d1_softwarereset~0 (
	.dataa(!\software_reset_request~q ),
	.datab(!\control[12]~q ),
	.datac(!\d1_softwarereset~q ),
	.datad(!\set_software_reset_bit~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d1_softwarereset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d1_softwarereset~0 .extended_lut = "off";
defparam \d1_softwarereset~0 .lut_mask = 64'h0A220A220A220A22;
defparam \d1_softwarereset~0 .shared_arith = "off";

dffeas d1_softwarereset(
	.clk(outclk_wire_0),
	.d(\d1_softwarereset~0_combout ),
	.asdata(vcc),
	.clrn(!system_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d1_softwarereset~q ),
	.prn(vcc));
defparam d1_softwarereset.is_wysiwyg = "true";
defparam d1_softwarereset.power_up = "low";

cyclonev_lcell_comb \software_reset_request~0 (
	.dataa(!\software_reset_request~q ),
	.datab(!\d1_softwarereset~q ),
	.datac(!\set_software_reset_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\software_reset_request~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \software_reset_request~0 .extended_lut = "off";
defparam \software_reset_request~0 .lut_mask = 64'h0202020202020202;
defparam \software_reset_request~0 .shared_arith = "off";

dffeas software_reset_request(
	.clk(outclk_wire_0),
	.d(\software_reset_request~0_combout ),
	.asdata(vcc),
	.clrn(!system_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\software_reset_request~q ),
	.prn(vcc));
defparam software_reset_request.is_wysiwyg = "true";
defparam software_reset_request.power_up = "low";

cyclonev_lcell_comb \reset_n~0 (
	.dataa(!\software_reset_request~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\reset_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \reset_n~0 .extended_lut = "off";
defparam \reset_n~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reset_n~0 .shared_arith = "off";

dffeas reset_n(
	.clk(outclk_wire_0),
	.d(\reset_n~0_combout ),
	.asdata(vcc),
	.clrn(!system_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_n~q ),
	.prn(vcc));
defparam reset_n.is_wysiwyg = "true";
defparam reset_n.power_up = "low";

dffeas \control[9] (
	.clk(outclk_wire_0),
	.d(in_data_reg_9),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[9]~q ),
	.prn(vcc));
defparam \control[9] .is_wysiwyg = "true";
defparam \control[9] .power_up = "low";

cyclonev_lcell_comb \Add1~125 (
	.dataa(!control_0),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[9]~q ),
	.datae(gnd),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~125_sumout ),
	.cout(\Add1~126 ),
	.shareout());
defparam \Add1~125 .extended_lut = "off";
defparam \Add1~125 .lut_mask = 64'h0000FF0000005500;
defparam \Add1~125 .shared_arith = "off";

cyclonev_lcell_comb \Add1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~121_sumout ),
	.cout(\Add1~122 ),
	.shareout());
defparam \Add1~121 .extended_lut = "off";
defparam \Add1~121 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~121 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!control_2),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[9]~q ),
	.datae(gnd),
	.dataf(!writeaddress_2),
	.datag(gnd),
	.cin(\Add1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000AA00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h0808080808080808;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_writeaddress~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writeaddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writeaddress~0 .extended_lut = "off";
defparam \p1_writeaddress~0 .lut_mask = 64'h0000000800000008;
defparam \p1_writeaddress~0 .shared_arith = "off";

cyclonev_lcell_comb \writeaddress[9]~0 (
	.dataa(!fifo_read),
	.datab(!\p1_writeaddress~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writeaddress[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writeaddress[9]~0 .extended_lut = "off";
defparam \writeaddress[9]~0 .lut_mask = 64'h7777777777777777;
defparam \writeaddress[9]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~37 .shared_arith = "off";

cyclonev_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout());
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~41 .shared_arith = "off";

cyclonev_lcell_comb \Add1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~45_sumout ),
	.cout(\Add1~46 ),
	.shareout());
defparam \Add1~45 .extended_lut = "off";
defparam \Add1~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~45 .shared_arith = "off";

cyclonev_lcell_comb \Add1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~49_sumout ),
	.cout(\Add1~50 ),
	.shareout());
defparam \Add1~49 .extended_lut = "off";
defparam \Add1~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~49 .shared_arith = "off";

cyclonev_lcell_comb \Add1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~53_sumout ),
	.cout(\Add1~54 ),
	.shareout());
defparam \Add1~53 .extended_lut = "off";
defparam \Add1~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~53 .shared_arith = "off";

cyclonev_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~57_sumout ),
	.cout(\Add1~58 ),
	.shareout());
defparam \Add1~57 .extended_lut = "off";
defparam \Add1~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~57 .shared_arith = "off";

cyclonev_lcell_comb \Add1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~61_sumout ),
	.cout(\Add1~62 ),
	.shareout());
defparam \Add1~61 .extended_lut = "off";
defparam \Add1~61 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~61 .shared_arith = "off";

cyclonev_lcell_comb \Add1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~65_sumout ),
	.cout(\Add1~66 ),
	.shareout());
defparam \Add1~65 .extended_lut = "off";
defparam \Add1~65 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~65 .shared_arith = "off";

cyclonev_lcell_comb \Add1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~69_sumout ),
	.cout(\Add1~70 ),
	.shareout());
defparam \Add1~69 .extended_lut = "off";
defparam \Add1~69 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~69 .shared_arith = "off";

cyclonev_lcell_comb \Add1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~73_sumout ),
	.cout(\Add1~74 ),
	.shareout());
defparam \Add1~73 .extended_lut = "off";
defparam \Add1~73 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~73 .shared_arith = "off";

cyclonev_lcell_comb \Add1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~77_sumout ),
	.cout(\Add1~78 ),
	.shareout());
defparam \Add1~77 .extended_lut = "off";
defparam \Add1~77 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~77 .shared_arith = "off";

cyclonev_lcell_comb \Add1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~81_sumout ),
	.cout(\Add1~82 ),
	.shareout());
defparam \Add1~81 .extended_lut = "off";
defparam \Add1~81 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~81 .shared_arith = "off";

cyclonev_lcell_comb \Add1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~85_sumout ),
	.cout(\Add1~86 ),
	.shareout());
defparam \Add1~85 .extended_lut = "off";
defparam \Add1~85 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~85 .shared_arith = "off";

cyclonev_lcell_comb \Add1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~89_sumout ),
	.cout(\Add1~90 ),
	.shareout());
defparam \Add1~89 .extended_lut = "off";
defparam \Add1~89 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~89 .shared_arith = "off";

cyclonev_lcell_comb \Add1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~93_sumout ),
	.cout(\Add1~94 ),
	.shareout());
defparam \Add1~93 .extended_lut = "off";
defparam \Add1~93 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~93 .shared_arith = "off";

cyclonev_lcell_comb \Add1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~97_sumout ),
	.cout(\Add1~98 ),
	.shareout());
defparam \Add1~97 .extended_lut = "off";
defparam \Add1~97 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~97 .shared_arith = "off";

cyclonev_lcell_comb \Add1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~101_sumout ),
	.cout(\Add1~102 ),
	.shareout());
defparam \Add1~101 .extended_lut = "off";
defparam \Add1~101 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~101 .shared_arith = "off";

cyclonev_lcell_comb \Add1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~105_sumout ),
	.cout(\Add1~106 ),
	.shareout());
defparam \Add1~105 .extended_lut = "off";
defparam \Add1~105 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~105 .shared_arith = "off";

cyclonev_lcell_comb \Add1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~109_sumout ),
	.cout(\Add1~110 ),
	.shareout());
defparam \Add1~109 .extended_lut = "off";
defparam \Add1~109 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~109 .shared_arith = "off";

cyclonev_lcell_comb \Add1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~113_sumout ),
	.cout(\Add1~114 ),
	.shareout());
defparam \Add1~113 .extended_lut = "off";
defparam \Add1~113 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~113 .shared_arith = "off";

cyclonev_lcell_comb \Add1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!writeaddress_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~117_sumout ),
	.cout(),
	.shareout());
defparam \Add1~117 .extended_lut = "off";
defparam \Add1~117 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~117 .shared_arith = "off";

dffeas \control[8] (
	.clk(outclk_wire_0),
	.d(in_data_reg_8),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[8]~q ),
	.prn(vcc));
defparam \control[8] .is_wysiwyg = "true";
defparam \control[8] .power_up = "low";

cyclonev_lcell_comb \Add0~61 (
	.dataa(!control_0),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[8]~q ),
	.datae(gnd),
	.dataf(!\readaddress[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0000005500;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~1 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~1 .extended_lut = "off";
defparam \Equal3~1 .lut_mask = 64'h4040404040404040;
defparam \Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_readaddress~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_readaddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_readaddress~0 .extended_lut = "off";
defparam \p1_readaddress~0 .lut_mask = 64'h0000000800000008;
defparam \p1_readaddress~0 .shared_arith = "off";

cyclonev_lcell_comb \readaddress[13]~0 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!\Equal3~1_combout ),
	.dataf(!read_latency_shift_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readaddress[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readaddress[13]~0 .extended_lut = "off";
defparam \readaddress[13]~0 .lut_mask = 64'h00000008FFFFFFFF;
defparam \readaddress[13]~0 .shared_arith = "off";

dffeas \readaddress[0] (
	.clk(outclk_wire_0),
	.d(\Add0~61_sumout ),
	.asdata(in_data_reg_0),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[0]~q ),
	.prn(vcc));
defparam \readaddress[0] .is_wysiwyg = "true";
defparam \readaddress[0] .power_up = "low";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~57 .shared_arith = "off";

dffeas \readaddress[1] (
	.clk(outclk_wire_0),
	.d(\Add0~57_sumout ),
	.asdata(in_data_reg_1),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[1]~q ),
	.prn(vcc));
defparam \readaddress[1] .is_wysiwyg = "true";
defparam \readaddress[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!control_2),
	.datab(gnd),
	.datac(gnd),
	.datad(!\control[8]~q ),
	.datae(gnd),
	.dataf(!readaddress_2),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF000000AA00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!readaddress_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \control[2]~0 (
	.dataa(!in_data_reg_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\control[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \control[2]~0 .extended_lut = "off";
defparam \control[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \control[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_0),
	.datad(!\writelength[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~113_sumout ),
	.cout(\Add3~114 ),
	.shareout(\Add3~115 ));
defparam \Add3~113 .extended_lut = "off";
defparam \Add3~113 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~113 .shared_arith = "on";

dffeas \writelength[30] (
	.clk(outclk_wire_0),
	.d(in_data_reg_30),
	.asdata(\Add3~1_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[30]~q ),
	.prn(vcc));
defparam \writelength[30] .is_wysiwyg = "true";
defparam \writelength[30] .power_up = "low";

cyclonev_lcell_comb \Add3~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~114 ),
	.sharein(\Add3~115 ),
	.combout(),
	.sumout(\Add3~117_sumout ),
	.cout(\Add3~118 ),
	.shareout(\Add3~119 ));
defparam \Add3~117 .extended_lut = "off";
defparam \Add3~117 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~117 .shared_arith = "on";

dffeas \writelength[1] (
	.clk(outclk_wire_0),
	.d(in_data_reg_1),
	.asdata(\Add3~117_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[1]~q ),
	.prn(vcc));
defparam \writelength[1] .is_wysiwyg = "true";
defparam \writelength[1] .power_up = "low";

cyclonev_lcell_comb \Add3~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!control_2),
	.datad(!\writelength[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~118 ),
	.sharein(\Add3~119 ),
	.combout(),
	.sumout(\Add3~121_sumout ),
	.cout(\Add3~122 ),
	.shareout(\Add3~123 ));
defparam \Add3~121 .extended_lut = "off";
defparam \Add3~121 .lut_mask = 64'h0000000F00000FF0;
defparam \Add3~121 .shared_arith = "on";

dffeas \writelength[2] (
	.clk(outclk_wire_0),
	.d(in_data_reg_2),
	.asdata(\Add3~121_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[2]~q ),
	.prn(vcc));
defparam \writelength[2] .is_wysiwyg = "true";
defparam \writelength[2] .power_up = "low";

cyclonev_lcell_comb \Add3~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~122 ),
	.sharein(\Add3~123 ),
	.combout(),
	.sumout(\Add3~125_sumout ),
	.cout(\Add3~126 ),
	.shareout(\Add3~127 ));
defparam \Add3~125 .extended_lut = "off";
defparam \Add3~125 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~125 .shared_arith = "on";

dffeas \writelength[3] (
	.clk(outclk_wire_0),
	.d(in_data_reg_3),
	.asdata(\Add3~125_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[3]~q ),
	.prn(vcc));
defparam \writelength[3] .is_wysiwyg = "true";
defparam \writelength[3] .power_up = "low";

cyclonev_lcell_comb \Add3~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~126 ),
	.sharein(\Add3~127 ),
	.combout(),
	.sumout(\Add3~49_sumout ),
	.cout(\Add3~50 ),
	.shareout(\Add3~51 ));
defparam \Add3~49 .extended_lut = "off";
defparam \Add3~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~49 .shared_arith = "on";

dffeas \writelength[4] (
	.clk(outclk_wire_0),
	.d(in_data_reg_4),
	.asdata(\Add3~49_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[4]~q ),
	.prn(vcc));
defparam \writelength[4] .is_wysiwyg = "true";
defparam \writelength[4] .power_up = "low";

cyclonev_lcell_comb \Add3~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~50 ),
	.sharein(\Add3~51 ),
	.combout(),
	.sumout(\Add3~53_sumout ),
	.cout(\Add3~54 ),
	.shareout(\Add3~55 ));
defparam \Add3~53 .extended_lut = "off";
defparam \Add3~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~53 .shared_arith = "on";

dffeas \writelength[5] (
	.clk(outclk_wire_0),
	.d(in_data_reg_5),
	.asdata(\Add3~53_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[5]~q ),
	.prn(vcc));
defparam \writelength[5] .is_wysiwyg = "true";
defparam \writelength[5] .power_up = "low";

cyclonev_lcell_comb \Add3~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~54 ),
	.sharein(\Add3~55 ),
	.combout(),
	.sumout(\Add3~57_sumout ),
	.cout(\Add3~58 ),
	.shareout(\Add3~59 ));
defparam \Add3~57 .extended_lut = "off";
defparam \Add3~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~57 .shared_arith = "on";

dffeas \writelength[6] (
	.clk(outclk_wire_0),
	.d(in_data_reg_6),
	.asdata(\Add3~57_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[6]~q ),
	.prn(vcc));
defparam \writelength[6] .is_wysiwyg = "true";
defparam \writelength[6] .power_up = "low";

cyclonev_lcell_comb \Add3~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~58 ),
	.sharein(\Add3~59 ),
	.combout(),
	.sumout(\Add3~61_sumout ),
	.cout(\Add3~62 ),
	.shareout(\Add3~63 ));
defparam \Add3~61 .extended_lut = "off";
defparam \Add3~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~61 .shared_arith = "on";

dffeas \writelength[7] (
	.clk(outclk_wire_0),
	.d(in_data_reg_7),
	.asdata(\Add3~61_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[7]~q ),
	.prn(vcc));
defparam \writelength[7] .is_wysiwyg = "true";
defparam \writelength[7] .power_up = "low";

cyclonev_lcell_comb \Add3~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~62 ),
	.sharein(\Add3~63 ),
	.combout(),
	.sumout(\Add3~65_sumout ),
	.cout(\Add3~66 ),
	.shareout(\Add3~67 ));
defparam \Add3~65 .extended_lut = "off";
defparam \Add3~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~65 .shared_arith = "on";

dffeas \writelength[8] (
	.clk(outclk_wire_0),
	.d(in_data_reg_8),
	.asdata(\Add3~65_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[8]~q ),
	.prn(vcc));
defparam \writelength[8] .is_wysiwyg = "true";
defparam \writelength[8] .power_up = "low";

cyclonev_lcell_comb \Add3~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~66 ),
	.sharein(\Add3~67 ),
	.combout(),
	.sumout(\Add3~69_sumout ),
	.cout(\Add3~70 ),
	.shareout(\Add3~71 ));
defparam \Add3~69 .extended_lut = "off";
defparam \Add3~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~69 .shared_arith = "on";

dffeas \writelength[9] (
	.clk(outclk_wire_0),
	.d(in_data_reg_9),
	.asdata(\Add3~69_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[9]~q ),
	.prn(vcc));
defparam \writelength[9] .is_wysiwyg = "true";
defparam \writelength[9] .power_up = "low";

cyclonev_lcell_comb \Add3~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~70 ),
	.sharein(\Add3~71 ),
	.combout(),
	.sumout(\Add3~93_sumout ),
	.cout(\Add3~94 ),
	.shareout(\Add3~95 ));
defparam \Add3~93 .extended_lut = "off";
defparam \Add3~93 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~93 .shared_arith = "on";

dffeas \writelength[10] (
	.clk(outclk_wire_0),
	.d(in_data_reg_10),
	.asdata(\Add3~93_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[10]~q ),
	.prn(vcc));
defparam \writelength[10] .is_wysiwyg = "true";
defparam \writelength[10] .power_up = "low";

cyclonev_lcell_comb \Add3~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~94 ),
	.sharein(\Add3~95 ),
	.combout(),
	.sumout(\Add3~97_sumout ),
	.cout(\Add3~98 ),
	.shareout(\Add3~99 ));
defparam \Add3~97 .extended_lut = "off";
defparam \Add3~97 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~97 .shared_arith = "on";

dffeas \writelength[11] (
	.clk(outclk_wire_0),
	.d(in_data_reg_11),
	.asdata(\Add3~97_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[11]~q ),
	.prn(vcc));
defparam \writelength[11] .is_wysiwyg = "true";
defparam \writelength[11] .power_up = "low";

cyclonev_lcell_comb \Add3~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~98 ),
	.sharein(\Add3~99 ),
	.combout(),
	.sumout(\Add3~101_sumout ),
	.cout(\Add3~102 ),
	.shareout(\Add3~103 ));
defparam \Add3~101 .extended_lut = "off";
defparam \Add3~101 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~101 .shared_arith = "on";

dffeas \writelength[12] (
	.clk(outclk_wire_0),
	.d(in_data_reg_12),
	.asdata(\Add3~101_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[12]~q ),
	.prn(vcc));
defparam \writelength[12] .is_wysiwyg = "true";
defparam \writelength[12] .power_up = "low";

cyclonev_lcell_comb \Add3~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~102 ),
	.sharein(\Add3~103 ),
	.combout(),
	.sumout(\Add3~105_sumout ),
	.cout(\Add3~106 ),
	.shareout(\Add3~107 ));
defparam \Add3~105 .extended_lut = "off";
defparam \Add3~105 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~105 .shared_arith = "on";

dffeas \writelength[13] (
	.clk(outclk_wire_0),
	.d(in_data_reg_13),
	.asdata(\Add3~105_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[13]~q ),
	.prn(vcc));
defparam \writelength[13] .is_wysiwyg = "true";
defparam \writelength[13] .power_up = "low";

cyclonev_lcell_comb \Add3~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~106 ),
	.sharein(\Add3~107 ),
	.combout(),
	.sumout(\Add3~109_sumout ),
	.cout(\Add3~110 ),
	.shareout(\Add3~111 ));
defparam \Add3~109 .extended_lut = "off";
defparam \Add3~109 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~109 .shared_arith = "on";

dffeas \writelength[14] (
	.clk(outclk_wire_0),
	.d(in_data_reg_14),
	.asdata(\Add3~109_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[14]~q ),
	.prn(vcc));
defparam \writelength[14] .is_wysiwyg = "true";
defparam \writelength[14] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~110 ),
	.sharein(\Add3~111 ),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout(\Add3~31 ));
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~29 .shared_arith = "on";

dffeas \writelength[15] (
	.clk(outclk_wire_0),
	.d(in_data_reg_15),
	.asdata(\Add3~29_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[15]~q ),
	.prn(vcc));
defparam \writelength[15] .is_wysiwyg = "true";
defparam \writelength[15] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(\Add3~31 ),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout(\Add3~35 ));
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~33 .shared_arith = "on";

dffeas \writelength[16] (
	.clk(outclk_wire_0),
	.d(in_data_reg_16),
	.asdata(\Add3~33_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[16]~q ),
	.prn(vcc));
defparam \writelength[16] .is_wysiwyg = "true";
defparam \writelength[16] .power_up = "low";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(\Add3~35 ),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout(\Add3~39 ));
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~37 .shared_arith = "on";

dffeas \writelength[17] (
	.clk(outclk_wire_0),
	.d(in_data_reg_17),
	.asdata(\Add3~37_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[17]~q ),
	.prn(vcc));
defparam \writelength[17] .is_wysiwyg = "true";
defparam \writelength[17] .power_up = "low";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(\Add3~39 ),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout(\Add3~43 ));
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~41 .shared_arith = "on";

dffeas \writelength[18] (
	.clk(outclk_wire_0),
	.d(in_data_reg_18),
	.asdata(\Add3~41_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[18]~q ),
	.prn(vcc));
defparam \writelength[18] .is_wysiwyg = "true";
defparam \writelength[18] .power_up = "low";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(\Add3~43 ),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout(\Add3~47 ));
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~45 .shared_arith = "on";

dffeas \writelength[19] (
	.clk(outclk_wire_0),
	.d(in_data_reg_19),
	.asdata(\Add3~45_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[19]~q ),
	.prn(vcc));
defparam \writelength[19] .is_wysiwyg = "true";
defparam \writelength[19] .power_up = "low";

cyclonev_lcell_comb \Add3~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(\Add3~47 ),
	.combout(),
	.sumout(\Add3~73_sumout ),
	.cout(\Add3~74 ),
	.shareout(\Add3~75 ));
defparam \Add3~73 .extended_lut = "off";
defparam \Add3~73 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~73 .shared_arith = "on";

dffeas \writelength[20] (
	.clk(outclk_wire_0),
	.d(in_data_reg_20),
	.asdata(\Add3~73_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[20]~q ),
	.prn(vcc));
defparam \writelength[20] .is_wysiwyg = "true";
defparam \writelength[20] .power_up = "low";

cyclonev_lcell_comb \Add3~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~74 ),
	.sharein(\Add3~75 ),
	.combout(),
	.sumout(\Add3~77_sumout ),
	.cout(\Add3~78 ),
	.shareout(\Add3~79 ));
defparam \Add3~77 .extended_lut = "off";
defparam \Add3~77 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~77 .shared_arith = "on";

dffeas \writelength[21] (
	.clk(outclk_wire_0),
	.d(in_data_reg_21),
	.asdata(\Add3~77_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[21]~q ),
	.prn(vcc));
defparam \writelength[21] .is_wysiwyg = "true";
defparam \writelength[21] .power_up = "low";

cyclonev_lcell_comb \Add3~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~78 ),
	.sharein(\Add3~79 ),
	.combout(),
	.sumout(\Add3~81_sumout ),
	.cout(\Add3~82 ),
	.shareout(\Add3~83 ));
defparam \Add3~81 .extended_lut = "off";
defparam \Add3~81 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~81 .shared_arith = "on";

dffeas \writelength[22] (
	.clk(outclk_wire_0),
	.d(in_data_reg_22),
	.asdata(\Add3~81_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[22]~q ),
	.prn(vcc));
defparam \writelength[22] .is_wysiwyg = "true";
defparam \writelength[22] .power_up = "low";

cyclonev_lcell_comb \Add3~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~82 ),
	.sharein(\Add3~83 ),
	.combout(),
	.sumout(\Add3~85_sumout ),
	.cout(\Add3~86 ),
	.shareout(\Add3~87 ));
defparam \Add3~85 .extended_lut = "off";
defparam \Add3~85 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~85 .shared_arith = "on";

dffeas \writelength[23] (
	.clk(outclk_wire_0),
	.d(in_data_reg_23),
	.asdata(\Add3~85_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[23]~q ),
	.prn(vcc));
defparam \writelength[23] .is_wysiwyg = "true";
defparam \writelength[23] .power_up = "low";

cyclonev_lcell_comb \Add3~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~86 ),
	.sharein(\Add3~87 ),
	.combout(),
	.sumout(\Add3~89_sumout ),
	.cout(\Add3~90 ),
	.shareout(\Add3~91 ));
defparam \Add3~89 .extended_lut = "off";
defparam \Add3~89 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~89 .shared_arith = "on";

dffeas \writelength[24] (
	.clk(outclk_wire_0),
	.d(in_data_reg_24),
	.asdata(\Add3~89_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[24]~q ),
	.prn(vcc));
defparam \writelength[24] .is_wysiwyg = "true";
defparam \writelength[24] .power_up = "low";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~90 ),
	.sharein(\Add3~91 ),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout(\Add3~11 ));
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~9 .shared_arith = "on";

dffeas \writelength[25] (
	.clk(outclk_wire_0),
	.d(in_data_reg_25),
	.asdata(\Add3~9_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[25]~q ),
	.prn(vcc));
defparam \writelength[25] .is_wysiwyg = "true";
defparam \writelength[25] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(\Add3~11 ),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout(\Add3~15 ));
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~13 .shared_arith = "on";

dffeas \writelength[26] (
	.clk(outclk_wire_0),
	.d(in_data_reg_26),
	.asdata(\Add3~13_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[26]~q ),
	.prn(vcc));
defparam \writelength[26] .is_wysiwyg = "true";
defparam \writelength[26] .power_up = "low";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(\Add3~15 ),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout(\Add3~19 ));
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~17 .shared_arith = "on";

dffeas \writelength[27] (
	.clk(outclk_wire_0),
	.d(in_data_reg_27),
	.asdata(\Add3~17_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[27]~q ),
	.prn(vcc));
defparam \writelength[27] .is_wysiwyg = "true";
defparam \writelength[27] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(\Add3~19 ),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout(\Add3~23 ));
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~21 .shared_arith = "on";

dffeas \writelength[28] (
	.clk(outclk_wire_0),
	.d(in_data_reg_28),
	.asdata(\Add3~21_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[28]~q ),
	.prn(vcc));
defparam \writelength[28] .is_wysiwyg = "true";
defparam \writelength[28] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(\Add3~23 ),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout(\Add3~27 ));
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~25 .shared_arith = "on";

dffeas \writelength[29] (
	.clk(outclk_wire_0),
	.d(in_data_reg_29),
	.asdata(\Add3~25_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[29]~q ),
	.prn(vcc));
defparam \writelength[29] .is_wysiwyg = "true";
defparam \writelength[29] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(\Add3~27 ),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout(\Add3~3 ));
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add3~1 .shared_arith = "on";

dffeas \writelength[31] (
	.clk(outclk_wire_0),
	.d(in_data_reg_31),
	.asdata(\Add3~5_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[31]~q ),
	.prn(vcc));
defparam \writelength[31] .is_wysiwyg = "true";
defparam \writelength[31] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\writelength[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(\Add3~3 ),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h000000000000FF00;
defparam \Add3~5 .shared_arith = "on";

cyclonev_lcell_comb \p1_writelength_eq_0~0 (
	.dataa(!\Add3~49_sumout ),
	.datab(!\Add3~53_sumout ),
	.datac(!\Add3~57_sumout ),
	.datad(!\Add3~61_sumout ),
	.datae(!\Add3~65_sumout ),
	.dataf(!\Add3~69_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~0 .extended_lut = "off";
defparam \p1_writelength_eq_0~0 .lut_mask = 64'h8000000000000000;
defparam \p1_writelength_eq_0~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~1 (
	.dataa(!\Add3~29_sumout ),
	.datab(!\Add3~33_sumout ),
	.datac(!\Add3~37_sumout ),
	.datad(!\Add3~41_sumout ),
	.datae(!\Add3~45_sumout ),
	.dataf(!\p1_writelength_eq_0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~1 .extended_lut = "off";
defparam \p1_writelength_eq_0~1 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~2 (
	.dataa(!\Add3~9_sumout ),
	.datab(!\Add3~13_sumout ),
	.datac(!\Add3~17_sumout ),
	.datad(!\Add3~21_sumout ),
	.datae(!\Add3~25_sumout ),
	.dataf(!\p1_writelength_eq_0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~2 .extended_lut = "off";
defparam \p1_writelength_eq_0~2 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~3 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!\Add3~113_sumout ),
	.datad(!\Add3~117_sumout ),
	.datae(!\Add3~121_sumout ),
	.dataf(!\Add3~125_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~3 .extended_lut = "off";
defparam \p1_writelength_eq_0~3 .lut_mask = 64'h1000000000000000;
defparam \p1_writelength_eq_0~3 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~4 (
	.dataa(!\Add3~93_sumout ),
	.datab(!\Add3~97_sumout ),
	.datac(!\Add3~101_sumout ),
	.datad(!\Add3~105_sumout ),
	.datae(!\Add3~109_sumout ),
	.dataf(!\p1_writelength_eq_0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~4 .extended_lut = "off";
defparam \p1_writelength_eq_0~4 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~4 .shared_arith = "off";

cyclonev_lcell_comb \p1_writelength_eq_0~5 (
	.dataa(!\Add3~73_sumout ),
	.datab(!\Add3~77_sumout ),
	.datac(!\Add3~81_sumout ),
	.datad(!\Add3~85_sumout ),
	.datae(!\Add3~89_sumout ),
	.dataf(!\p1_writelength_eq_0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_writelength_eq_0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_writelength_eq_0~5 .extended_lut = "off";
defparam \p1_writelength_eq_0~5 .lut_mask = 64'h0000000080000000;
defparam \p1_writelength_eq_0~5 .shared_arith = "off";

cyclonev_lcell_comb \writelength_eq_0~0 (
	.dataa(!\writelength_eq_0~q ),
	.datab(!\Add3~1_sumout ),
	.datac(!\Add3~5_sumout ),
	.datad(!\p1_writelength_eq_0~2_combout ),
	.datae(!\p1_writelength_eq_0~5_combout ),
	.dataf(!\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writelength_eq_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writelength_eq_0~0 .extended_lut = "off";
defparam \writelength_eq_0~0 .lut_mask = 64'hFFFFFFFF55555515;
defparam \writelength_eq_0~0 .shared_arith = "off";

dffeas writelength_eq_0(
	.clk(outclk_wire_0),
	.d(\writelength_eq_0~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writelength_eq_0~q ),
	.prn(vcc));
defparam writelength_eq_0.is_wysiwyg = "true";
defparam writelength_eq_0.power_up = "low";

cyclonev_lcell_comb \writelength[8]~0 (
	.dataa(!fifo_read),
	.datab(!\writelength_eq_0~q ),
	.datac(!\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\writelength[8]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \writelength[8]~0 .extended_lut = "off";
defparam \writelength[8]~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \writelength[8]~0 .shared_arith = "off";

dffeas \writelength[0] (
	.clk(outclk_wire_0),
	.d(in_data_reg_0),
	.asdata(\Add3~113_sumout ),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\the_Computer_System_dma_2_read_data_mux|length_write~combout ),
	.ena(\writelength[8]~0_combout ),
	.q(\writelength[0]~q ),
	.prn(vcc));
defparam \writelength[0] .is_wysiwyg = "true";
defparam \writelength[0] .power_up = "low";

cyclonev_lcell_comb \Equal3~2 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~2 .extended_lut = "off";
defparam \Equal3~2 .lut_mask = 64'h0404040404040404;
defparam \Equal3~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[0]~0 (
	.dataa(!writeaddress_0),
	.datab(!\Equal3~0_combout ),
	.datac(!\readaddress[0]~q ),
	.datad(!\Equal3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[0]~0 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[0]~0 .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~3 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~3 .extended_lut = "off";
defparam \Equal3~3 .lut_mask = 64'h0202020202020202;
defparam \Equal3~3 .shared_arith = "off";

dffeas \control[3] (
	.clk(outclk_wire_0),
	.d(in_data_reg_3),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[3]~q ),
	.prn(vcc));
defparam \control[3] .is_wysiwyg = "true";
defparam \control[3] .power_up = "low";

cyclonev_lcell_comb \control[7]~1 (
	.dataa(!in_data_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\control[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \control[7]~1 .extended_lut = "off";
defparam \control[7]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \control[7]~1 .shared_arith = "off";

dffeas \control[7] (
	.clk(outclk_wire_0),
	.d(\control[7]~1_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[7]~q ),
	.prn(vcc));
defparam \control[7] .is_wysiwyg = "true";
defparam \control[7] .power_up = "low";

cyclonev_lcell_comb \p1_done_write~0 (
	.dataa(!\control[7]~q ),
	.datab(!\writelength_eq_0~q ),
	.datac(!\Add3~1_sumout ),
	.datad(!\Add3~5_sumout ),
	.datae(!\p1_writelength_eq_0~2_combout ),
	.dataf(!\p1_writelength_eq_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_done_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_done_write~0 .extended_lut = "off";
defparam \p1_done_write~0 .lut_mask = 64'h888888888888A888;
defparam \p1_done_write~0 .shared_arith = "off";

dffeas done_write(
	.clk(outclk_wire_0),
	.d(\p1_done_write~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\done_write~q ),
	.prn(vcc));
defparam done_write.is_wysiwyg = "true";
defparam done_write.power_up = "low";

cyclonev_lcell_comb done_transaction(
	.dataa(!\control[3]~q ),
	.datab(!\done_write~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\done_transaction~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam done_transaction.extended_lut = "off";
defparam done_transaction.lut_mask = 64'h1111111111111111;
defparam done_transaction.shared_arith = "off";

dffeas d1_done_transaction(
	.clk(outclk_wire_0),
	.d(\done_transaction~combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d1_done_transaction~q ),
	.prn(vcc));
defparam d1_done_transaction.is_wysiwyg = "true";
defparam d1_done_transaction.power_up = "low";

cyclonev_lcell_comb flush_fifo(
	.dataa(!\control[3]~q ),
	.datab(!\done_write~q ),
	.datac(!\d1_done_transaction~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\flush_fifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam flush_fifo.extended_lut = "off";
defparam flush_fifo.lut_mask = 64'h1010101010101010;
defparam flush_fifo.shared_arith = "off";

cyclonev_lcell_comb \p1_readaddress~1 (
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_readaddress~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_readaddress~1 .extended_lut = "off";
defparam \p1_readaddress~1 .lut_mask = 64'h0008000800080008;
defparam \p1_readaddress~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata~1 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata~1 .extended_lut = "off";
defparam \p1_dma_ctl_readdata~1 .lut_mask = 64'h8080808080808080;
defparam \p1_dma_ctl_readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \done~0 (
	.dataa(!\flush_fifo~combout ),
	.datab(!\p1_readaddress~1_combout ),
	.datac(!\done~q ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \done~0 .extended_lut = "off";
defparam \done~0 .lut_mask = 64'h5F4C5F4C5F4C5F4C;
defparam \done~0 .shared_arith = "off";

dffeas done(
	.clk(outclk_wire_0),
	.d(\done~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\done~q ),
	.prn(vcc));
defparam done.is_wysiwyg = "true";
defparam done.power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[0]~2 (
	.dataa(!control_0),
	.datab(!\Equal3~3_combout ),
	.datac(!\done~q ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[0]~2 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[0]~2 .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[0] (
	.dataa(!\writelength[0]~q ),
	.datab(!\Equal3~2_combout ),
	.datac(!\p1_dma_ctl_readdata[0]~0_combout ),
	.datad(!\p1_dma_ctl_readdata[0]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[0] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[0] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \p1_dma_ctl_readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[1]~3 (
	.dataa(!writeaddress_1),
	.datab(!\Equal3~0_combout ),
	.datac(!\readaddress[1]~q ),
	.datad(!\Equal3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[1]~3 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[1]~3 .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[1]~3 .shared_arith = "off";

dffeas \control[1] (
	.clk(outclk_wire_0),
	.d(in_data_reg_1),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[1]~q ),
	.prn(vcc));
defparam \control[1] .is_wysiwyg = "true";
defparam \control[1] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[1]~4 (
	.dataa(!\control[3]~q ),
	.datab(!\done_write~q ),
	.datac(!\Equal3~3_combout ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(!\control[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[1]~4 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[1]~4 .lut_mask = 64'h00440F4F00440F4F;
defparam \p1_dma_ctl_readdata[1]~4 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[1] (
	.dataa(!\writelength[1]~q ),
	.datab(!\Equal3~2_combout ),
	.datac(!\p1_dma_ctl_readdata[1]~3_combout ),
	.datad(!\p1_dma_ctl_readdata[1]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[1] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[1] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \p1_dma_ctl_readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[2]~43 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_2),
	.datad(!\writelength[2]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!control_2),
	.datag(!readaddress_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[2]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[2]~43 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[2]~43 .lut_mask = 64'h02024C6E0202082A;
defparam \p1_dma_ctl_readdata[2]~43 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[3]~39 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_3),
	.datad(!\writelength[3]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\control[3]~q ),
	.datag(!readaddress_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[3]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[3]~39 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[3]~39 .lut_mask = 64'h0202082A02024C6E;
defparam \p1_dma_ctl_readdata[3]~39 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[4]~5 (
	.dataa(!writeaddress_4),
	.datab(!readaddress_4),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[4]~5 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[4]~5 .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[4]~5 .shared_arith = "off";

dffeas \control[4] (
	.clk(outclk_wire_0),
	.d(in_data_reg_4),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[4]~q ),
	.prn(vcc));
defparam \control[4] .is_wysiwyg = "true";
defparam \control[4] .power_up = "low";

cyclonev_lcell_comb \len~0 (
	.dataa(!\flush_fifo~combout ),
	.datab(!\p1_readaddress~1_combout ),
	.datac(!\writelength_eq_0~q ),
	.datad(!\p1_dma_ctl_readdata~1_combout ),
	.datae(!\len~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\len~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \len~0 .extended_lut = "off";
defparam \len~0 .lut_mask = 64'h5040FFCC5040FFCC;
defparam \len~0 .shared_arith = "off";

dffeas len(
	.clk(outclk_wire_0),
	.d(\len~0_combout ),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\len~q ),
	.prn(vcc));
defparam len.is_wysiwyg = "true";
defparam len.power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[4]~6 (
	.dataa(!\Equal3~3_combout ),
	.datab(!\p1_dma_ctl_readdata~1_combout ),
	.datac(!\control[4]~q ),
	.datad(!\len~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[4]~6 .extended_lut = "off";
defparam \p1_dma_ctl_readdata[4]~6 .lut_mask = 64'h0537053705370537;
defparam \p1_dma_ctl_readdata[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[4] (
	.dataa(!\writelength[4]~q ),
	.datab(!\Equal3~2_combout ),
	.datac(!\p1_dma_ctl_readdata[4]~5_combout ),
	.datad(!\p1_dma_ctl_readdata[4]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[4] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[4] .lut_mask = 64'h1FFF1FFF1FFF1FFF;
defparam \p1_dma_ctl_readdata[4] .shared_arith = "off";

dffeas \control[5] (
	.clk(outclk_wire_0),
	.d(in_data_reg_5),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[5]~q ),
	.prn(vcc));
defparam \control[5] .is_wysiwyg = "true";
defparam \control[5] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[5]~35 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_5),
	.datad(!\control[5]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[5]~q ),
	.datag(!readaddress_5),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[5]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[5]~35 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[5]~35 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[5]~35 .shared_arith = "off";

dffeas \control[6] (
	.clk(outclk_wire_0),
	.d(in_data_reg_6),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[6]~q ),
	.prn(vcc));
defparam \control[6] .is_wysiwyg = "true";
defparam \control[6] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[6]~31 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_6),
	.datad(!\control[6]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[6]~q ),
	.datag(!readaddress_6),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[6]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[6]~31 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[6]~31 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[6]~31 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[7]~27 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_7),
	.datad(!\writelength[7]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\control[7]~q ),
	.datag(!readaddress_7),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[7]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[7]~27 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[7]~27 .lut_mask = 64'h02024C6E0202082A;
defparam \p1_dma_ctl_readdata[7]~27 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[8]~23 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_8),
	.datad(!\writelength[8]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\control[8]~q ),
	.datag(!readaddress_8),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[8]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[8]~23 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[8]~23 .lut_mask = 64'h0202082A02024C6E;
defparam \p1_dma_ctl_readdata[8]~23 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[9]~19 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_9),
	.datad(!\writelength[9]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\control[9]~q ),
	.datag(!readaddress_9),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[9]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[9]~19 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[9]~19 .lut_mask = 64'h0202082A02024C6E;
defparam \p1_dma_ctl_readdata[9]~19 .shared_arith = "off";

dffeas \control[10] (
	.clk(outclk_wire_0),
	.d(in_data_reg_10),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[10]~q ),
	.prn(vcc));
defparam \control[10] .is_wysiwyg = "true";
defparam \control[10] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[10]~15 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_10),
	.datad(!\control[10]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[10]~q ),
	.datag(!readaddress_10),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[10]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[10]~15 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[10]~15 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[10]~15 .shared_arith = "off";

dffeas \control[11] (
	.clk(outclk_wire_0),
	.d(in_data_reg_11),
	.asdata(vcc),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p1_control~0_combout ),
	.q(\control[11]~q ),
	.prn(vcc));
defparam \control[11] .is_wysiwyg = "true";
defparam \control[11] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[11]~11 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_11),
	.datad(!\control[11]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[11]~q ),
	.datag(!readaddress_11),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[11]~11 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[11]~11 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[11]~11 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[12]~7 (
	.dataa(!int_nxt_addr_reg_dly_4),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!writeaddress_12),
	.datad(!\control[12]~q ),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[12]~q ),
	.datag(!readaddress_12),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[12]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[12]~7 .extended_lut = "on";
defparam \p1_dma_ctl_readdata[12]~7 .lut_mask = 64'h0202084C02022A6E;
defparam \p1_dma_ctl_readdata[12]~7 .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[13] (
	.dataa(!writeaddress_13),
	.datab(!readaddress_13),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[13]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[13] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[13] .lut_mask = 64'h0300500003005F00;
defparam \p1_dma_ctl_readdata[13] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[14] (
	.dataa(!writeaddress_14),
	.datab(!readaddress_14),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[14] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[14] .lut_mask = 64'h0300500003005F00;
defparam \p1_dma_ctl_readdata[14] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[15] (
	.dataa(!writeaddress_15),
	.datab(!readaddress_15),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(!int_nxt_addr_reg_dly_3),
	.dataf(!\writelength[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[15] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[15] .lut_mask = 64'h0300500003005F00;
defparam \p1_dma_ctl_readdata[15] .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~65 .shared_arith = "off";

dffeas \readaddress[16] (
	.clk(outclk_wire_0),
	.d(\Add0~65_sumout ),
	.asdata(in_data_reg_16),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[16]~q ),
	.prn(vcc));
defparam \readaddress[16] .is_wysiwyg = "true";
defparam \readaddress[16] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[16] (
	.dataa(!writeaddress_16),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[16]~q ),
	.dataf(!\readaddress[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[16] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[16] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[16] .shared_arith = "off";

cyclonev_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~69 .shared_arith = "off";

dffeas \readaddress[17] (
	.clk(outclk_wire_0),
	.d(\Add0~69_sumout ),
	.asdata(in_data_reg_17),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[17]~q ),
	.prn(vcc));
defparam \readaddress[17] .is_wysiwyg = "true";
defparam \readaddress[17] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[17] (
	.dataa(!writeaddress_17),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[17]~q ),
	.dataf(!\readaddress[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[17] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[17] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[17] .shared_arith = "off";

cyclonev_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~73 .shared_arith = "off";

dffeas \readaddress[18] (
	.clk(outclk_wire_0),
	.d(\Add0~73_sumout ),
	.asdata(in_data_reg_18),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[18]~q ),
	.prn(vcc));
defparam \readaddress[18] .is_wysiwyg = "true";
defparam \readaddress[18] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[18] (
	.dataa(!writeaddress_18),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[18]~q ),
	.dataf(!\readaddress[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[18] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[18] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[18] .shared_arith = "off";

cyclonev_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~77 .shared_arith = "off";

dffeas \readaddress[19] (
	.clk(outclk_wire_0),
	.d(\Add0~77_sumout ),
	.asdata(in_data_reg_19),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[19]~q ),
	.prn(vcc));
defparam \readaddress[19] .is_wysiwyg = "true";
defparam \readaddress[19] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[19] (
	.dataa(!writeaddress_19),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[19]~q ),
	.dataf(!\readaddress[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[19] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[19] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[19] .shared_arith = "off";

cyclonev_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~81 .shared_arith = "off";

dffeas \readaddress[20] (
	.clk(outclk_wire_0),
	.d(\Add0~81_sumout ),
	.asdata(in_data_reg_20),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[20]~q ),
	.prn(vcc));
defparam \readaddress[20] .is_wysiwyg = "true";
defparam \readaddress[20] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[20] (
	.dataa(!writeaddress_20),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[20]~q ),
	.dataf(!\readaddress[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[20] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[20] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[20] .shared_arith = "off";

cyclonev_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~85 .shared_arith = "off";

dffeas \readaddress[21] (
	.clk(outclk_wire_0),
	.d(\Add0~85_sumout ),
	.asdata(in_data_reg_21),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[21]~q ),
	.prn(vcc));
defparam \readaddress[21] .is_wysiwyg = "true";
defparam \readaddress[21] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[21] (
	.dataa(!writeaddress_21),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[21]~q ),
	.dataf(!\readaddress[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[21] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[21] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[21] .shared_arith = "off";

cyclonev_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~89 .shared_arith = "off";

dffeas \readaddress[22] (
	.clk(outclk_wire_0),
	.d(\Add0~89_sumout ),
	.asdata(in_data_reg_22),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[22]~q ),
	.prn(vcc));
defparam \readaddress[22] .is_wysiwyg = "true";
defparam \readaddress[22] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[22] (
	.dataa(!writeaddress_22),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[22]~q ),
	.dataf(!\readaddress[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[22] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[22] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[22] .shared_arith = "off";

cyclonev_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~93 .shared_arith = "off";

dffeas \readaddress[23] (
	.clk(outclk_wire_0),
	.d(\Add0~93_sumout ),
	.asdata(in_data_reg_23),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[23]~q ),
	.prn(vcc));
defparam \readaddress[23] .is_wysiwyg = "true";
defparam \readaddress[23] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[23] (
	.dataa(!writeaddress_23),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[23]~q ),
	.dataf(!\readaddress[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[23] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[23] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[23] .shared_arith = "off";

cyclonev_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~97 .shared_arith = "off";

dffeas \readaddress[24] (
	.clk(outclk_wire_0),
	.d(\Add0~97_sumout ),
	.asdata(in_data_reg_24),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[24]~q ),
	.prn(vcc));
defparam \readaddress[24] .is_wysiwyg = "true";
defparam \readaddress[24] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[24] (
	.dataa(!writeaddress_24),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[24]~q ),
	.dataf(!\readaddress[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[24] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[24] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[24] .shared_arith = "off";

cyclonev_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~101 .shared_arith = "off";

dffeas \readaddress[25] (
	.clk(outclk_wire_0),
	.d(\Add0~101_sumout ),
	.asdata(in_data_reg_25),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[25]~q ),
	.prn(vcc));
defparam \readaddress[25] .is_wysiwyg = "true";
defparam \readaddress[25] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[25] (
	.dataa(!writeaddress_25),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[25]~q ),
	.dataf(!\readaddress[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[25] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[25] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[25] .shared_arith = "off";

cyclonev_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~105 .shared_arith = "off";

dffeas \readaddress[26] (
	.clk(outclk_wire_0),
	.d(\Add0~105_sumout ),
	.asdata(in_data_reg_26),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[26]~q ),
	.prn(vcc));
defparam \readaddress[26] .is_wysiwyg = "true";
defparam \readaddress[26] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[26] (
	.dataa(!writeaddress_26),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[26]~q ),
	.dataf(!\readaddress[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[26] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[26] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[26] .shared_arith = "off";

cyclonev_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\readaddress[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~109 .shared_arith = "off";

dffeas \readaddress[27] (
	.clk(outclk_wire_0),
	.d(\Add0~109_sumout ),
	.asdata(in_data_reg_27),
	.clrn(\reset_n~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\p1_readaddress~0_combout ),
	.ena(\readaddress[13]~0_combout ),
	.q(\readaddress[27]~q ),
	.prn(vcc));
defparam \readaddress[27] .is_wysiwyg = "true";
defparam \readaddress[27] .power_up = "low";

cyclonev_lcell_comb \p1_dma_ctl_readdata[27] (
	.dataa(!writeaddress_27),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\writelength[27]~q ),
	.dataf(!\readaddress[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[27] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[27] .lut_mask = 64'h0040007030403070;
defparam \p1_dma_ctl_readdata[27] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[28] (
	.dataa(!writeaddress_28),
	.datab(!\Equal3~0_combout ),
	.datac(!\writelength[28]~q ),
	.datad(!\Equal3~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[28] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[28] .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[28] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[29] (
	.dataa(!writeaddress_29),
	.datab(!\Equal3~0_combout ),
	.datac(!\writelength[29]~q ),
	.datad(!\Equal3~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[29] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[29] .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[29] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[30] (
	.dataa(!writeaddress_30),
	.datab(!\Equal3~0_combout ),
	.datac(!\writelength[30]~q ),
	.datad(!\Equal3~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[30] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[30] .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[30] .shared_arith = "off";

cyclonev_lcell_comb \p1_dma_ctl_readdata[31] (
	.dataa(!writeaddress_31),
	.datab(!\Equal3~0_combout ),
	.datac(!\writelength[31]~q ),
	.datad(!\Equal3~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_dma_ctl_readdata[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_dma_ctl_readdata[31] .extended_lut = "off";
defparam \p1_dma_ctl_readdata[31] .lut_mask = 64'h111F111F111F111F;
defparam \p1_dma_ctl_readdata[31] .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_2_fifo_module (
	outclk_wire_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	fifo_empty1,
	src_valid,
	last_write_collision1,
	last_write_data_0,
	last_write_data_1,
	last_write_data_2,
	last_write_data_3,
	last_write_data_4,
	last_write_data_5,
	last_write_data_6,
	last_write_data_7,
	last_write_data_8,
	last_write_data_9,
	last_write_data_10,
	last_write_data_11,
	last_write_data_12,
	last_write_data_13,
	last_write_data_14,
	last_write_data_15,
	last_write_data_16,
	last_write_data_17,
	last_write_data_18,
	last_write_data_19,
	last_write_data_20,
	last_write_data_21,
	last_write_data_22,
	last_write_data_23,
	last_write_data_24,
	last_write_data_25,
	last_write_data_26,
	last_write_data_27,
	last_write_data_28,
	last_write_data_29,
	last_write_data_30,
	last_write_data_31,
	fifo_read,
	write_cp_ready,
	flush_fifo,
	src0_valid,
	reset_n,
	l1_w16_n0_mux_dataout,
	fifo_wr_data_0,
	l1_w17_n0_mux_dataout,
	fifo_wr_data_1,
	l1_w18_n0_mux_dataout,
	fifo_wr_data_2,
	l1_w19_n0_mux_dataout,
	fifo_wr_data_3,
	l1_w20_n0_mux_dataout,
	fifo_wr_data_4,
	l1_w21_n0_mux_dataout,
	fifo_wr_data_5,
	l1_w22_n0_mux_dataout,
	fifo_wr_data_6,
	l1_w23_n0_mux_dataout,
	fifo_wr_data_7,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout,
	read_latency_shift_reg,
	p1_fifo_full)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	fifo_empty1;
input 	src_valid;
output 	last_write_collision1;
output 	last_write_data_0;
output 	last_write_data_1;
output 	last_write_data_2;
output 	last_write_data_3;
output 	last_write_data_4;
output 	last_write_data_5;
output 	last_write_data_6;
output 	last_write_data_7;
output 	last_write_data_8;
output 	last_write_data_9;
output 	last_write_data_10;
output 	last_write_data_11;
output 	last_write_data_12;
output 	last_write_data_13;
output 	last_write_data_14;
output 	last_write_data_15;
output 	last_write_data_16;
output 	last_write_data_17;
output 	last_write_data_18;
output 	last_write_data_19;
output 	last_write_data_20;
output 	last_write_data_21;
output 	last_write_data_22;
output 	last_write_data_23;
output 	last_write_data_24;
output 	last_write_data_25;
output 	last_write_data_26;
output 	last_write_data_27;
output 	last_write_data_28;
output 	last_write_data_29;
output 	last_write_data_30;
output 	last_write_data_31;
input 	fifo_read;
input 	write_cp_ready;
input 	flush_fifo;
input 	src0_valid;
input 	reset_n;
input 	l1_w16_n0_mux_dataout;
input 	fifo_wr_data_0;
input 	l1_w17_n0_mux_dataout;
input 	fifo_wr_data_1;
input 	l1_w18_n0_mux_dataout;
input 	fifo_wr_data_2;
input 	l1_w19_n0_mux_dataout;
input 	fifo_wr_data_3;
input 	l1_w20_n0_mux_dataout;
input 	fifo_wr_data_4;
input 	l1_w21_n0_mux_dataout;
input 	fifo_wr_data_5;
input 	l1_w22_n0_mux_dataout;
input 	fifo_wr_data_6;
input 	l1_w23_n0_mux_dataout;
input 	fifo_wr_data_7;
input 	l1_w8_n0_mux_dataout;
input 	l1_w9_n0_mux_dataout;
input 	l1_w10_n0_mux_dataout;
input 	l1_w11_n0_mux_dataout;
input 	l1_w12_n0_mux_dataout;
input 	l1_w13_n0_mux_dataout;
input 	l1_w14_n0_mux_dataout;
input 	l1_w15_n0_mux_dataout;
input 	l1_w24_n0_mux_dataout;
input 	l1_w25_n0_mux_dataout;
input 	l1_w26_n0_mux_dataout;
input 	l1_w27_n0_mux_dataout;
input 	l1_w28_n0_mux_dataout;
input 	l1_w29_n0_mux_dataout;
input 	l1_w30_n0_mux_dataout;
input 	l1_w31_n0_mux_dataout;
input 	read_latency_shift_reg;
output 	p1_fifo_full;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wraddress~3_combout ;
wire \wraddress[1]~1_combout ;
wire \wraddress[0]~q ;
wire \wraddress~4_combout ;
wire \wraddress[1]~q ;
wire \wraddress~5_combout ;
wire \wraddress[2]~q ;
wire \wraddress~0_combout ;
wire \wraddress[3]~q ;
wire \rdaddress[0]~1_combout ;
wire \rdaddress_reg[0]~q ;
wire \rdaddress[1]~2_combout ;
wire \rdaddress_reg[1]~q ;
wire \Add1~1_combout ;
wire \rdaddress[2]~3_combout ;
wire \rdaddress_reg[2]~q ;
wire \Add1~0_combout ;
wire \rdaddress[3]~4_combout ;
wire \rdaddress_reg[3]~q ;
wire \wraddress~2_combout ;
wire \wraddress[4]~q ;
wire \Add1~2_combout ;
wire \rdaddress[4]~0_combout ;
wire \rdaddress_reg[4]~q ;
wire \p1_fifo_empty~0_combout ;
wire \p1_fifo_empty~1_combout ;
wire \p1_fifo_empty~2_combout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \write_collision~0_combout ;
wire \write_collision~combout ;
wire \last_write_collision~0_combout ;
wire \estimated_wraddress~4_combout ;
wire \estimated_wraddress[1]~1_combout ;
wire \estimated_wraddress[0]~q ;
wire \estimated_wraddress~5_combout ;
wire \estimated_wraddress[1]~q ;
wire \estimated_wraddress~2_combout ;
wire \estimated_wraddress[2]~q ;
wire \estimated_wraddress~3_combout ;
wire \estimated_wraddress[3]~q ;
wire \estimated_wraddress~0_combout ;
wire \estimated_wraddress[4]~q ;
wire \fifo_full~q ;
wire \p1_fifo_full~0_combout ;
wire \p1_fifo_full~1_combout ;
wire \p1_fifo_full~2_combout ;


Computer_System_Computer_System_dma_2_fifo_module_fifo_ram_module Computer_System_dma_2_fifo_module_fifo_ram(
	.outclk_wire_0(outclk_wire_0),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.src0_valid(src0_valid),
	.wraddress_3(\wraddress[3]~q ),
	.wraddress_4(\wraddress[4]~q ),
	.wraddress_0(\wraddress[0]~q ),
	.wraddress_1(\wraddress[1]~q ),
	.wraddress_2(\wraddress[2]~q ),
	.rdaddress_4(\rdaddress[4]~0_combout ),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout),
	.fifo_wr_data_0(fifo_wr_data_0),
	.rdaddress_0(\rdaddress[0]~1_combout ),
	.rdaddress_1(\rdaddress[1]~2_combout ),
	.rdaddress_2(\rdaddress[2]~3_combout ),
	.rdaddress_3(\rdaddress[3]~4_combout ),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout),
	.fifo_wr_data_1(fifo_wr_data_1),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout),
	.fifo_wr_data_2(fifo_wr_data_2),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout),
	.fifo_wr_data_3(fifo_wr_data_3),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout),
	.fifo_wr_data_4(fifo_wr_data_4),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout),
	.fifo_wr_data_5(fifo_wr_data_5),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout),
	.fifo_wr_data_6(fifo_wr_data_6),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout),
	.fifo_wr_data_7(fifo_wr_data_7),
	.l1_w8_n0_mux_dataout(l1_w8_n0_mux_dataout),
	.l1_w9_n0_mux_dataout(l1_w9_n0_mux_dataout),
	.l1_w10_n0_mux_dataout(l1_w10_n0_mux_dataout),
	.l1_w11_n0_mux_dataout(l1_w11_n0_mux_dataout),
	.l1_w12_n0_mux_dataout(l1_w12_n0_mux_dataout),
	.l1_w13_n0_mux_dataout(l1_w13_n0_mux_dataout),
	.l1_w14_n0_mux_dataout(l1_w14_n0_mux_dataout),
	.l1_w15_n0_mux_dataout(l1_w15_n0_mux_dataout),
	.l1_w24_n0_mux_dataout(l1_w24_n0_mux_dataout),
	.l1_w25_n0_mux_dataout(l1_w25_n0_mux_dataout),
	.l1_w26_n0_mux_dataout(l1_w26_n0_mux_dataout),
	.l1_w27_n0_mux_dataout(l1_w27_n0_mux_dataout),
	.l1_w28_n0_mux_dataout(l1_w28_n0_mux_dataout),
	.l1_w29_n0_mux_dataout(l1_w29_n0_mux_dataout),
	.l1_w30_n0_mux_dataout(l1_w30_n0_mux_dataout),
	.l1_w31_n0_mux_dataout(l1_w31_n0_mux_dataout));

dffeas fifo_empty(
	.clk(outclk_wire_0),
	.d(\p1_fifo_empty~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_empty1),
	.prn(vcc));
defparam fifo_empty.is_wysiwyg = "true";
defparam fifo_empty.power_up = "low";

dffeas last_write_collision(
	.clk(outclk_wire_0),
	.d(\last_write_collision~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_write_collision1),
	.prn(vcc));
defparam last_write_collision.is_wysiwyg = "true";
defparam last_write_collision.power_up = "low";

dffeas \last_write_data[0] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_0),
	.prn(vcc));
defparam \last_write_data[0] .is_wysiwyg = "true";
defparam \last_write_data[0] .power_up = "low";

dffeas \last_write_data[1] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_1),
	.prn(vcc));
defparam \last_write_data[1] .is_wysiwyg = "true";
defparam \last_write_data[1] .power_up = "low";

dffeas \last_write_data[2] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_2),
	.prn(vcc));
defparam \last_write_data[2] .is_wysiwyg = "true";
defparam \last_write_data[2] .power_up = "low";

dffeas \last_write_data[3] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_3),
	.prn(vcc));
defparam \last_write_data[3] .is_wysiwyg = "true";
defparam \last_write_data[3] .power_up = "low";

dffeas \last_write_data[4] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_4),
	.prn(vcc));
defparam \last_write_data[4] .is_wysiwyg = "true";
defparam \last_write_data[4] .power_up = "low";

dffeas \last_write_data[5] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_5),
	.prn(vcc));
defparam \last_write_data[5] .is_wysiwyg = "true";
defparam \last_write_data[5] .power_up = "low";

dffeas \last_write_data[6] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_6),
	.prn(vcc));
defparam \last_write_data[6] .is_wysiwyg = "true";
defparam \last_write_data[6] .power_up = "low";

dffeas \last_write_data[7] (
	.clk(outclk_wire_0),
	.d(fifo_wr_data_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_7),
	.prn(vcc));
defparam \last_write_data[7] .is_wysiwyg = "true";
defparam \last_write_data[7] .power_up = "low";

dffeas \last_write_data[8] (
	.clk(outclk_wire_0),
	.d(l1_w8_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_8),
	.prn(vcc));
defparam \last_write_data[8] .is_wysiwyg = "true";
defparam \last_write_data[8] .power_up = "low";

dffeas \last_write_data[9] (
	.clk(outclk_wire_0),
	.d(l1_w9_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_9),
	.prn(vcc));
defparam \last_write_data[9] .is_wysiwyg = "true";
defparam \last_write_data[9] .power_up = "low";

dffeas \last_write_data[10] (
	.clk(outclk_wire_0),
	.d(l1_w10_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_10),
	.prn(vcc));
defparam \last_write_data[10] .is_wysiwyg = "true";
defparam \last_write_data[10] .power_up = "low";

dffeas \last_write_data[11] (
	.clk(outclk_wire_0),
	.d(l1_w11_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_11),
	.prn(vcc));
defparam \last_write_data[11] .is_wysiwyg = "true";
defparam \last_write_data[11] .power_up = "low";

dffeas \last_write_data[12] (
	.clk(outclk_wire_0),
	.d(l1_w12_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_12),
	.prn(vcc));
defparam \last_write_data[12] .is_wysiwyg = "true";
defparam \last_write_data[12] .power_up = "low";

dffeas \last_write_data[13] (
	.clk(outclk_wire_0),
	.d(l1_w13_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_13),
	.prn(vcc));
defparam \last_write_data[13] .is_wysiwyg = "true";
defparam \last_write_data[13] .power_up = "low";

dffeas \last_write_data[14] (
	.clk(outclk_wire_0),
	.d(l1_w14_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_14),
	.prn(vcc));
defparam \last_write_data[14] .is_wysiwyg = "true";
defparam \last_write_data[14] .power_up = "low";

dffeas \last_write_data[15] (
	.clk(outclk_wire_0),
	.d(l1_w15_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_15),
	.prn(vcc));
defparam \last_write_data[15] .is_wysiwyg = "true";
defparam \last_write_data[15] .power_up = "low";

dffeas \last_write_data[16] (
	.clk(outclk_wire_0),
	.d(l1_w16_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_16),
	.prn(vcc));
defparam \last_write_data[16] .is_wysiwyg = "true";
defparam \last_write_data[16] .power_up = "low";

dffeas \last_write_data[17] (
	.clk(outclk_wire_0),
	.d(l1_w17_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_17),
	.prn(vcc));
defparam \last_write_data[17] .is_wysiwyg = "true";
defparam \last_write_data[17] .power_up = "low";

dffeas \last_write_data[18] (
	.clk(outclk_wire_0),
	.d(l1_w18_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_18),
	.prn(vcc));
defparam \last_write_data[18] .is_wysiwyg = "true";
defparam \last_write_data[18] .power_up = "low";

dffeas \last_write_data[19] (
	.clk(outclk_wire_0),
	.d(l1_w19_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_19),
	.prn(vcc));
defparam \last_write_data[19] .is_wysiwyg = "true";
defparam \last_write_data[19] .power_up = "low";

dffeas \last_write_data[20] (
	.clk(outclk_wire_0),
	.d(l1_w20_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_20),
	.prn(vcc));
defparam \last_write_data[20] .is_wysiwyg = "true";
defparam \last_write_data[20] .power_up = "low";

dffeas \last_write_data[21] (
	.clk(outclk_wire_0),
	.d(l1_w21_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_21),
	.prn(vcc));
defparam \last_write_data[21] .is_wysiwyg = "true";
defparam \last_write_data[21] .power_up = "low";

dffeas \last_write_data[22] (
	.clk(outclk_wire_0),
	.d(l1_w22_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_22),
	.prn(vcc));
defparam \last_write_data[22] .is_wysiwyg = "true";
defparam \last_write_data[22] .power_up = "low";

dffeas \last_write_data[23] (
	.clk(outclk_wire_0),
	.d(l1_w23_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_23),
	.prn(vcc));
defparam \last_write_data[23] .is_wysiwyg = "true";
defparam \last_write_data[23] .power_up = "low";

dffeas \last_write_data[24] (
	.clk(outclk_wire_0),
	.d(l1_w24_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_24),
	.prn(vcc));
defparam \last_write_data[24] .is_wysiwyg = "true";
defparam \last_write_data[24] .power_up = "low";

dffeas \last_write_data[25] (
	.clk(outclk_wire_0),
	.d(l1_w25_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_25),
	.prn(vcc));
defparam \last_write_data[25] .is_wysiwyg = "true";
defparam \last_write_data[25] .power_up = "low";

dffeas \last_write_data[26] (
	.clk(outclk_wire_0),
	.d(l1_w26_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_26),
	.prn(vcc));
defparam \last_write_data[26] .is_wysiwyg = "true";
defparam \last_write_data[26] .power_up = "low";

dffeas \last_write_data[27] (
	.clk(outclk_wire_0),
	.d(l1_w27_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_27),
	.prn(vcc));
defparam \last_write_data[27] .is_wysiwyg = "true";
defparam \last_write_data[27] .power_up = "low";

dffeas \last_write_data[28] (
	.clk(outclk_wire_0),
	.d(l1_w28_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_28),
	.prn(vcc));
defparam \last_write_data[28] .is_wysiwyg = "true";
defparam \last_write_data[28] .power_up = "low";

dffeas \last_write_data[29] (
	.clk(outclk_wire_0),
	.d(l1_w29_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_29),
	.prn(vcc));
defparam \last_write_data[29] .is_wysiwyg = "true";
defparam \last_write_data[29] .power_up = "low";

dffeas \last_write_data[30] (
	.clk(outclk_wire_0),
	.d(l1_w30_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_30),
	.prn(vcc));
defparam \last_write_data[30] .is_wysiwyg = "true";
defparam \last_write_data[30] .power_up = "low";

dffeas \last_write_data[31] (
	.clk(outclk_wire_0),
	.d(l1_w31_n0_mux_dataout),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_collision~combout ),
	.q(last_write_data_31),
	.prn(vcc));
defparam \last_write_data[31] .is_wysiwyg = "true";
defparam \last_write_data[31] .power_up = "low";

cyclonev_lcell_comb \p1_fifo_full~3 (
	.dataa(!flush_fifo),
	.datab(!\rdaddress[4]~0_combout ),
	.datac(!\estimated_wraddress[4]~q ),
	.datad(!\p1_fifo_full~0_combout ),
	.datae(!\p1_fifo_full~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(p1_fifo_full),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~3 .extended_lut = "off";
defparam \p1_fifo_full~3 .lut_mask = 64'h00AA28AA00AA28AA;
defparam \p1_fifo_full~3 .shared_arith = "off";

cyclonev_lcell_comb \wraddress~3 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~3 .extended_lut = "off";
defparam \wraddress~3 .lut_mask = 64'h8888888888888888;
defparam \wraddress~3 .shared_arith = "off";

cyclonev_lcell_comb \wraddress[1]~1 (
	.dataa(!flush_fifo),
	.datab(!src0_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress[1]~1 .extended_lut = "off";
defparam \wraddress[1]~1 .lut_mask = 64'h7777777777777777;
defparam \wraddress[1]~1 .shared_arith = "off";

dffeas \wraddress[0] (
	.clk(outclk_wire_0),
	.d(\wraddress~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[1]~1_combout ),
	.q(\wraddress[0]~q ),
	.prn(vcc));
defparam \wraddress[0] .is_wysiwyg = "true";
defparam \wraddress[0] .power_up = "low";

cyclonev_lcell_comb \wraddress~4 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~4 .extended_lut = "off";
defparam \wraddress~4 .lut_mask = 64'h8282828282828282;
defparam \wraddress~4 .shared_arith = "off";

dffeas \wraddress[1] (
	.clk(outclk_wire_0),
	.d(\wraddress~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[1]~1_combout ),
	.q(\wraddress[1]~q ),
	.prn(vcc));
defparam \wraddress[1] .is_wysiwyg = "true";
defparam \wraddress[1] .power_up = "low";

cyclonev_lcell_comb \wraddress~5 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\wraddress[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~5 .extended_lut = "off";
defparam \wraddress~5 .lut_mask = 64'h802A802A802A802A;
defparam \wraddress~5 .shared_arith = "off";

dffeas \wraddress[2] (
	.clk(outclk_wire_0),
	.d(\wraddress~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[1]~1_combout ),
	.q(\wraddress[2]~q ),
	.prn(vcc));
defparam \wraddress[2] .is_wysiwyg = "true";
defparam \wraddress[2] .power_up = "low";

cyclonev_lcell_comb \wraddress~0 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\wraddress[2]~q ),
	.datae(!\wraddress[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~0 .extended_lut = "off";
defparam \wraddress~0 .lut_mask = 64'h80002AAA80002AAA;
defparam \wraddress~0 .shared_arith = "off";

dffeas \wraddress[3] (
	.clk(outclk_wire_0),
	.d(\wraddress~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[1]~1_combout ),
	.q(\wraddress[3]~q ),
	.prn(vcc));
defparam \wraddress[3] .is_wysiwyg = "true";
defparam \wraddress[3] .power_up = "low";

cyclonev_lcell_comb \rdaddress[0]~1 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\rdaddress_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[0]~1 .extended_lut = "off";
defparam \rdaddress[0]~1 .lut_mask = 64'h10E010E010E010E0;
defparam \rdaddress[0]~1 .shared_arith = "off";

dffeas \rdaddress_reg[0] (
	.clk(outclk_wire_0),
	.d(\rdaddress[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[0]~q ),
	.prn(vcc));
defparam \rdaddress_reg[0] .is_wysiwyg = "true";
defparam \rdaddress_reg[0] .power_up = "low";

cyclonev_lcell_comb \rdaddress[1]~2 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\rdaddress_reg[0]~q ),
	.datae(!\rdaddress_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[1]~2 .extended_lut = "off";
defparam \rdaddress[1]~2 .lut_mask = 64'h1000E0F01000E0F0;
defparam \rdaddress[1]~2 .shared_arith = "off";

dffeas \rdaddress_reg[1] (
	.clk(outclk_wire_0),
	.d(\rdaddress[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[1]~q ),
	.prn(vcc));
defparam \rdaddress_reg[1] .is_wysiwyg = "true";
defparam \rdaddress_reg[1] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\rdaddress_reg[0]~q ),
	.datab(!\rdaddress_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h8888888888888888;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \rdaddress[2]~3 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\rdaddress_reg[2]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[2]~3 .extended_lut = "off";
defparam \rdaddress[2]~3 .lut_mask = 64'h00F010E000F010E0;
defparam \rdaddress[2]~3 .shared_arith = "off";

dffeas \rdaddress_reg[2] (
	.clk(outclk_wire_0),
	.d(\rdaddress[2]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[2]~q ),
	.prn(vcc));
defparam \rdaddress_reg[2] .is_wysiwyg = "true";
defparam \rdaddress_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\rdaddress_reg[0]~q ),
	.datab(!\rdaddress_reg[1]~q ),
	.datac(!\rdaddress_reg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8080808080808080;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \rdaddress[3]~4 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\rdaddress_reg[3]~q ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[3]~4 .extended_lut = "off";
defparam \rdaddress[3]~4 .lut_mask = 64'h00F010E000F010E0;
defparam \rdaddress[3]~4 .shared_arith = "off";

dffeas \rdaddress_reg[3] (
	.clk(outclk_wire_0),
	.d(\rdaddress[3]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[3]~q ),
	.prn(vcc));
defparam \rdaddress_reg[3] .is_wysiwyg = "true";
defparam \rdaddress_reg[3] .power_up = "low";

cyclonev_lcell_comb \wraddress~2 (
	.dataa(!flush_fifo),
	.datab(!\wraddress[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\wraddress[2]~q ),
	.datae(!\wraddress[3]~q ),
	.dataf(!\wraddress[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wraddress~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wraddress~2 .extended_lut = "off";
defparam \wraddress~2 .lut_mask = 64'h800000002AAAAAAA;
defparam \wraddress~2 .shared_arith = "off";

dffeas \wraddress[4] (
	.clk(outclk_wire_0),
	.d(\wraddress~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wraddress[1]~1_combout ),
	.q(\wraddress[4]~q ),
	.prn(vcc));
defparam \wraddress[4] .is_wysiwyg = "true";
defparam \wraddress[4] .power_up = "low";

cyclonev_lcell_comb \Add1~2 (
	.dataa(!\rdaddress_reg[0]~q ),
	.datab(!\rdaddress_reg[1]~q ),
	.datac(!\rdaddress_reg[2]~q ),
	.datad(!\rdaddress_reg[3]~q ),
	.datae(!\rdaddress_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~2 .extended_lut = "off";
defparam \Add1~2 .lut_mask = 64'h7FFF80007FFF8000;
defparam \Add1~2 .shared_arith = "off";

cyclonev_lcell_comb \rdaddress[4]~0 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\rdaddress_reg[4]~q ),
	.datae(!\Add1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdaddress[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdaddress[4]~0 .extended_lut = "off";
defparam \rdaddress[4]~0 .lut_mask = 64'h10F000E010F000E0;
defparam \rdaddress[4]~0 .shared_arith = "off";

dffeas \rdaddress_reg[4] (
	.clk(outclk_wire_0),
	.d(\rdaddress[4]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdaddress_reg[4]~q ),
	.prn(vcc));
defparam \rdaddress_reg[4] .is_wysiwyg = "true";
defparam \rdaddress_reg[4] .power_up = "low";

cyclonev_lcell_comb \p1_fifo_empty~0 (
	.dataa(!\wraddress[0]~q ),
	.datab(!\rdaddress_reg[0]~q ),
	.datac(!\wraddress[1]~q ),
	.datad(!\rdaddress_reg[1]~q ),
	.datae(!\wraddress[2]~q ),
	.dataf(!\rdaddress_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~0 .extended_lut = "off";
defparam \p1_fifo_empty~0 .lut_mask = 64'h2042040004002042;
defparam \p1_fifo_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_empty~1 (
	.dataa(!\wraddress[3]~q ),
	.datab(!\rdaddress_reg[3]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\wraddress[4]~q ),
	.datae(!\rdaddress_reg[4]~q ),
	.dataf(!\p1_fifo_empty~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~1 .extended_lut = "off";
defparam \p1_fifo_empty~1 .lut_mask = 64'h0000000092040492;
defparam \p1_fifo_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_empty~2 (
	.dataa(!fifo_empty1),
	.datab(!fifo_read),
	.datac(!flush_fifo),
	.datad(!src0_valid),
	.datae(!\p1_fifo_empty~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_empty~2 .extended_lut = "off";
defparam \p1_fifo_empty~2 .lut_mask = 64'h50F040F050F040F0;
defparam \p1_fifo_empty~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\rdaddress_reg[0]~q ),
	.datae(!\wraddress[1]~q ),
	.dataf(!\rdaddress_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h1000EFFFE0F01F0F;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\wraddress[2]~q ),
	.datae(!\rdaddress_reg[2]~q ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h00FFF00F10EFE01F;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~2 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!\wraddress[3]~q ),
	.datae(!\rdaddress_reg[3]~q ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~2 .extended_lut = "off";
defparam \Equal2~2 .lut_mask = 64'h00FFF00F10EFE01F;
defparam \Equal2~2 .shared_arith = "off";

cyclonev_lcell_comb \write_collision~0 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!flush_fifo),
	.datad(!src0_valid),
	.datae(!\wraddress[0]~q ),
	.dataf(!\rdaddress_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_collision~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_collision~0 .extended_lut = "off";
defparam \write_collision~0 .lut_mask = 64'h00EF0010001F00E0;
defparam \write_collision~0 .shared_arith = "off";

cyclonev_lcell_comb write_collision(
	.dataa(!\wraddress[4]~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\Equal2~1_combout ),
	.datad(!\Equal2~2_combout ),
	.datae(!\rdaddress[4]~0_combout ),
	.dataf(!\write_collision~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_collision~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam write_collision.extended_lut = "off";
defparam write_collision.lut_mask = 64'h0000000080004000;
defparam write_collision.shared_arith = "off";

cyclonev_lcell_comb \last_write_collision~0 (
	.dataa(!last_write_collision1),
	.datab(!fifo_read),
	.datac(!\write_collision~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_write_collision~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_write_collision~0 .extended_lut = "off";
defparam \last_write_collision~0 .lut_mask = 64'h4F4F4F4F4F4F4F4F;
defparam \last_write_collision~0 .shared_arith = "off";

cyclonev_lcell_comb \estimated_wraddress~4 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~4 .extended_lut = "off";
defparam \estimated_wraddress~4 .lut_mask = 64'h8888888888888888;
defparam \estimated_wraddress~4 .shared_arith = "off";

cyclonev_lcell_comb \estimated_wraddress[1]~1 (
	.dataa(!flush_fifo),
	.datab(!read_latency_shift_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress[1]~1 .extended_lut = "off";
defparam \estimated_wraddress[1]~1 .lut_mask = 64'h7777777777777777;
defparam \estimated_wraddress[1]~1 .shared_arith = "off";

dffeas \estimated_wraddress[0] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[1]~1_combout ),
	.q(\estimated_wraddress[0]~q ),
	.prn(vcc));
defparam \estimated_wraddress[0] .is_wysiwyg = "true";
defparam \estimated_wraddress[0] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~5 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~5 .extended_lut = "off";
defparam \estimated_wraddress~5 .lut_mask = 64'h2828282828282828;
defparam \estimated_wraddress~5 .shared_arith = "off";

dffeas \estimated_wraddress[1] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[1]~1_combout ),
	.q(\estimated_wraddress[1]~q ),
	.prn(vcc));
defparam \estimated_wraddress[1] .is_wysiwyg = "true";
defparam \estimated_wraddress[1] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~2 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\estimated_wraddress[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~2 .extended_lut = "off";
defparam \estimated_wraddress~2 .lut_mask = 64'h02A802A802A802A8;
defparam \estimated_wraddress~2 .shared_arith = "off";

dffeas \estimated_wraddress[2] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[1]~1_combout ),
	.q(\estimated_wraddress[2]~q ),
	.prn(vcc));
defparam \estimated_wraddress[2] .is_wysiwyg = "true";
defparam \estimated_wraddress[2] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~3 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\estimated_wraddress[2]~q ),
	.datae(!\estimated_wraddress[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~3 .extended_lut = "off";
defparam \estimated_wraddress~3 .lut_mask = 64'h0002AAA80002AAA8;
defparam \estimated_wraddress~3 .shared_arith = "off";

dffeas \estimated_wraddress[3] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[1]~1_combout ),
	.q(\estimated_wraddress[3]~q ),
	.prn(vcc));
defparam \estimated_wraddress[3] .is_wysiwyg = "true";
defparam \estimated_wraddress[3] .power_up = "low";

cyclonev_lcell_comb \estimated_wraddress~0 (
	.dataa(!flush_fifo),
	.datab(!\estimated_wraddress[0]~q ),
	.datac(!\estimated_wraddress[1]~q ),
	.datad(!\estimated_wraddress[2]~q ),
	.datae(!\estimated_wraddress[3]~q ),
	.dataf(!\estimated_wraddress[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\estimated_wraddress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \estimated_wraddress~0 .extended_lut = "off";
defparam \estimated_wraddress~0 .lut_mask = 64'h00000002AAAAAAA8;
defparam \estimated_wraddress~0 .shared_arith = "off";

dffeas \estimated_wraddress[4] (
	.clk(outclk_wire_0),
	.d(\estimated_wraddress~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\estimated_wraddress[1]~1_combout ),
	.q(\estimated_wraddress[4]~q ),
	.prn(vcc));
defparam \estimated_wraddress[4] .is_wysiwyg = "true";
defparam \estimated_wraddress[4] .power_up = "low";

dffeas fifo_full(
	.clk(outclk_wire_0),
	.d(p1_fifo_full),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_full~q ),
	.prn(vcc));
defparam fifo_full.is_wysiwyg = "true";
defparam fifo_full.power_up = "low";

cyclonev_lcell_comb \p1_fifo_full~0 (
	.dataa(!fifo_read),
	.datab(!src0_valid),
	.datac(!\fifo_full~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~0 .extended_lut = "off";
defparam \p1_fifo_full~0 .lut_mask = 64'h0B0B0B0B0B0B0B0B;
defparam \p1_fifo_full~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_full~1 (
	.dataa(!\rdaddress[0]~1_combout ),
	.datab(!\rdaddress[1]~2_combout ),
	.datac(!read_latency_shift_reg),
	.datad(!\estimated_wraddress[0]~q ),
	.datae(!\estimated_wraddress[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~1 .extended_lut = "off";
defparam \p1_fifo_full~1 .lut_mask = 64'h0102040801020408;
defparam \p1_fifo_full~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_fifo_full~2 (
	.dataa(!\rdaddress[2]~3_combout ),
	.datab(!\rdaddress[3]~4_combout ),
	.datac(!\estimated_wraddress[2]~q ),
	.datad(!\estimated_wraddress[3]~q ),
	.datae(!\p1_fifo_full~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_fifo_full~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_fifo_full~2 .extended_lut = "off";
defparam \p1_fifo_full~2 .lut_mask = 64'h0000124800001248;
defparam \p1_fifo_full~2 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_2_fifo_module_fifo_ram_module (
	outclk_wire_0,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	src0_valid,
	wraddress_3,
	wraddress_4,
	wraddress_0,
	wraddress_1,
	wraddress_2,
	rdaddress_4,
	l1_w16_n0_mux_dataout,
	fifo_wr_data_0,
	rdaddress_0,
	rdaddress_1,
	rdaddress_2,
	rdaddress_3,
	l1_w17_n0_mux_dataout,
	fifo_wr_data_1,
	l1_w18_n0_mux_dataout,
	fifo_wr_data_2,
	l1_w19_n0_mux_dataout,
	fifo_wr_data_3,
	l1_w20_n0_mux_dataout,
	fifo_wr_data_4,
	l1_w21_n0_mux_dataout,
	fifo_wr_data_5,
	l1_w22_n0_mux_dataout,
	fifo_wr_data_6,
	l1_w23_n0_mux_dataout,
	fifo_wr_data_7,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	src0_valid;
input 	wraddress_3;
input 	wraddress_4;
input 	wraddress_0;
input 	wraddress_1;
input 	wraddress_2;
input 	rdaddress_4;
input 	l1_w16_n0_mux_dataout;
input 	fifo_wr_data_0;
input 	rdaddress_0;
input 	rdaddress_1;
input 	rdaddress_2;
input 	rdaddress_3;
input 	l1_w17_n0_mux_dataout;
input 	fifo_wr_data_1;
input 	l1_w18_n0_mux_dataout;
input 	fifo_wr_data_2;
input 	l1_w19_n0_mux_dataout;
input 	fifo_wr_data_3;
input 	l1_w20_n0_mux_dataout;
input 	fifo_wr_data_4;
input 	l1_w21_n0_mux_dataout;
input 	fifo_wr_data_5;
input 	l1_w22_n0_mux_dataout;
input 	fifo_wr_data_6;
input 	l1_w23_n0_mux_dataout;
input 	fifo_wr_data_7;
input 	l1_w8_n0_mux_dataout;
input 	l1_w9_n0_mux_dataout;
input 	l1_w10_n0_mux_dataout;
input 	l1_w11_n0_mux_dataout;
input 	l1_w12_n0_mux_dataout;
input 	l1_w13_n0_mux_dataout;
input 	l1_w14_n0_mux_dataout;
input 	l1_w15_n0_mux_dataout;
input 	l1_w24_n0_mux_dataout;
input 	l1_w25_n0_mux_dataout;
input 	l1_w26_n0_mux_dataout;
input 	l1_w27_n0_mux_dataout;
input 	l1_w28_n0_mux_dataout;
input 	l1_w29_n0_mux_dataout;
input 	l1_w30_n0_mux_dataout;
input 	l1_w31_n0_mux_dataout;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_lpm_ram_dp_2 lpm_ram_dp_component(
	.wrclock(outclk_wire_0),
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren(src0_valid),
	.wraddress({wraddress_4,wraddress_3,wraddress_2,wraddress_1,wraddress_0}),
	.rdaddress({rdaddress_4,rdaddress_3,rdaddress_2,rdaddress_1,rdaddress_0}),
	.data({l1_w31_n0_mux_dataout,l1_w30_n0_mux_dataout,l1_w29_n0_mux_dataout,l1_w28_n0_mux_dataout,l1_w27_n0_mux_dataout,l1_w26_n0_mux_dataout,l1_w25_n0_mux_dataout,l1_w24_n0_mux_dataout,l1_w23_n0_mux_dataout,l1_w22_n0_mux_dataout,l1_w21_n0_mux_dataout,l1_w20_n0_mux_dataout,
l1_w19_n0_mux_dataout,l1_w18_n0_mux_dataout,l1_w17_n0_mux_dataout,l1_w16_n0_mux_dataout,l1_w15_n0_mux_dataout,l1_w14_n0_mux_dataout,l1_w13_n0_mux_dataout,l1_w12_n0_mux_dataout,l1_w11_n0_mux_dataout,l1_w10_n0_mux_dataout,l1_w9_n0_mux_dataout,l1_w8_n0_mux_dataout,
fifo_wr_data_7,fifo_wr_data_6,fifo_wr_data_5,fifo_wr_data_4,fifo_wr_data_3,fifo_wr_data_2,fifo_wr_data_1,fifo_wr_data_0}));

endmodule

module Computer_System_lpm_ram_dp_2 (
	wrclock,
	q,
	wren,
	wraddress,
	rdaddress,
	data)/* synthesis synthesis_greybox=0 */;
input 	wrclock;
output 	[31:0] q;
input 	wren;
input 	[4:0] wraddress;
input 	[4:0] rdaddress;
input 	[31:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdpram_2 sram(
	.inclock(wrclock),
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren(wren),
	.wraddress({wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.rdaddress({rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module Computer_System_altdpram_2 (
	inclock,
	q,
	wren,
	wraddress,
	rdaddress,
	data)/* synthesis synthesis_greybox=0 */;
input 	inclock;
output 	[31:0] q;
input 	wren;
input 	[4:0] wraddress;
input 	[4:0] rdaddress;
input 	[31:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altsyncram_2 ram_block(
	.clock0(inclock),
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren_a(wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,wraddress[4],wraddress[3],wraddress[2],wraddress[1],wraddress[0]}),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rdaddress[4],rdaddress[3],rdaddress[2],rdaddress[1],rdaddress[0]}),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module Computer_System_altsyncram_2 (
	clock0,
	q_b,
	wren_a,
	address_a,
	address_b,
	data_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
output 	[31:0] q_b;
input 	wren_a;
input 	[13:0] address_a;
input 	[13:0] address_b;
input 	[31:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altsyncram_1j02_1 auto_generated(
	.clock0(clock0),
	.clock1(clock0),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}));

endmodule

module Computer_System_altsyncram_1j02_1 (
	clock0,
	clock1,
	q_b,
	wren_a,
	address_a,
	address_b,
	data_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
input 	clock1;
output 	[31:0] q_b;
input 	wren_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	[31:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.clk1_input_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.clk1_input_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.clk1_input_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.clk1_input_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.clk1_input_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.clk1_input_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.clk1_input_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.clk1_input_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.clk1_input_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.clk1_input_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.clk1_input_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.clk1_input_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.clk1_input_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.clk1_input_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.clk1_input_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.clk1_input_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Computer_System_dma_2:dma_2|Computer_System_dma_2_fifo_module:the_Computer_System_dma_2_fifo_module|Computer_System_dma_2_fifo_module_fifo_ram_module:Computer_System_dma_2_fifo_module_fifo_ram|lpm_ram_dp:lpm_ram_dp_component|altdpram:sram|altsyncram:ram_block|altsyncram_1j02:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module Computer_System_Computer_System_dma_2_mem_read (
	clk,
	hold_waitrequest,
	saved_grant_0,
	mem_used_1,
	control_3,
	reset_n,
	read_select1,
	read_latency_shift_reg,
	control_7,
	p1_done_write,
	p1_done_read,
	p1_fifo_full)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	hold_waitrequest;
input 	saved_grant_0;
input 	mem_used_1;
input 	control_3;
input 	reset_n;
output 	read_select1;
input 	read_latency_shift_reg;
input 	control_7;
input 	p1_done_write;
input 	p1_done_read;
input 	p1_fifo_full;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \p1_read_select~0_combout ;
wire \Computer_System_dma_2_mem_read_idle~0_combout ;
wire \Computer_System_dma_2_mem_read_idle~4_combout ;
wire \Computer_System_dma_2_mem_read_idle~q ;
wire \Computer_System_dma_2_mem_read_access~0_combout ;
wire \p1_read_select~1_combout ;


dffeas read_select(
	.clk(clk),
	.d(\p1_read_select~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_select1),
	.prn(vcc));
defparam read_select.is_wysiwyg = "true";
defparam read_select.power_up = "low";

cyclonev_lcell_comb \p1_read_select~0 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!read_select1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_read_select~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_read_select~0 .extended_lut = "off";
defparam \p1_read_select~0 .lut_mask = 64'h00EF00EF00EF00EF;
defparam \p1_read_select~0 .shared_arith = "off";

cyclonev_lcell_comb \Computer_System_dma_2_mem_read_idle~0 (
	.dataa(!p1_fifo_full),
	.datab(!p1_done_read),
	.datac(!read_latency_shift_reg),
	.datad(!p1_done_write),
	.datae(!\Computer_System_dma_2_mem_read_idle~q ),
	.dataf(!control_7),
	.datag(!control_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_2_mem_read_idle~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_2_mem_read_idle~0 .extended_lut = "on";
defparam \Computer_System_dma_2_mem_read_idle~0 .lut_mask = 64'hFDFF0D0FF5F50505;
defparam \Computer_System_dma_2_mem_read_idle~0 .shared_arith = "off";

cyclonev_lcell_comb \Computer_System_dma_2_mem_read_idle~4 (
	.dataa(!\Computer_System_dma_2_mem_read_idle~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_2_mem_read_idle~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_2_mem_read_idle~4 .extended_lut = "off";
defparam \Computer_System_dma_2_mem_read_idle~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Computer_System_dma_2_mem_read_idle~4 .shared_arith = "off";

dffeas Computer_System_dma_2_mem_read_idle(
	.clk(clk),
	.d(\Computer_System_dma_2_mem_read_idle~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\Computer_System_dma_2_mem_read_idle~q ),
	.prn(vcc));
defparam Computer_System_dma_2_mem_read_idle.is_wysiwyg = "true";
defparam Computer_System_dma_2_mem_read_idle.power_up = "low";

cyclonev_lcell_comb \Computer_System_dma_2_mem_read_access~0 (
	.dataa(!control_3),
	.datab(!read_select1),
	.datac(!\Computer_System_dma_2_mem_read_idle~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Computer_System_dma_2_mem_read_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Computer_System_dma_2_mem_read_access~0 .extended_lut = "off";
defparam \Computer_System_dma_2_mem_read_access~0 .lut_mask = 64'h8C8C8C8C8C8C8C8C;
defparam \Computer_System_dma_2_mem_read_access~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_read_select~1 (
	.dataa(!control_7),
	.datab(!p1_done_write),
	.datac(!\p1_read_select~0_combout ),
	.datad(!\Computer_System_dma_2_mem_read_access~0_combout ),
	.datae(!p1_done_read),
	.dataf(!p1_fifo_full),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_read_select~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_read_select~1 .extended_lut = "off";
defparam \p1_read_select~1 .lut_mask = 64'h5F0FDF0F0F0F0F0F;
defparam \p1_read_select~1 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_2_mem_write (
	f2h_AWREADY_0,
	f2h_WREADY_0,
	address_taken,
	mem_used_7,
	src_valid,
	data_taken,
	fifo_read)/* synthesis synthesis_greybox=0 */;
input 	f2h_AWREADY_0;
input 	f2h_WREADY_0;
input 	address_taken;
input 	mem_used_7;
input 	src_valid;
input 	data_taken;
output 	fifo_read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \fifo_read~0 (
	.dataa(!f2h_AWREADY_0),
	.datab(!f2h_WREADY_0),
	.datac(!address_taken),
	.datad(!mem_used_7),
	.datae(!src_valid),
	.dataf(!data_taken),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_read),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_read~0 .extended_lut = "off";
defparam \fifo_read~0 .lut_mask = 64'h0000130300005757;
defparam \fifo_read~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_dma_2_read_data_mux (
	ram_block1a32,
	ram_block1a0,
	ram_block1a33,
	ram_block1a1,
	ram_block1a34,
	ram_block1a2,
	ram_block1a35,
	ram_block1a3,
	ram_block1a36,
	ram_block1a4,
	ram_block1a37,
	ram_block1a5,
	ram_block1a38,
	ram_block1a6,
	ram_block1a39,
	ram_block1a7,
	ram_block1a40,
	ram_block1a8,
	ram_block1a41,
	ram_block1a9,
	ram_block1a42,
	ram_block1a10,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a59,
	ram_block1a27,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	clk,
	readaddress_0,
	readaddress_1,
	control_2,
	control_0,
	WideOr0,
	wait_latency_counter_1,
	src0_valid,
	reset_n,
	in_data_reg_59,
	mem,
	in_data_reg_3,
	address_reg_a_0,
	l1_w16_n0_mux_dataout,
	fifo_wr_data_0,
	p1_control,
	l1_w17_n0_mux_dataout,
	fifo_wr_data_1,
	l1_w18_n0_mux_dataout,
	fifo_wr_data_2,
	l1_w19_n0_mux_dataout,
	fifo_wr_data_3,
	l1_w20_n0_mux_dataout,
	fifo_wr_data_4,
	l1_w21_n0_mux_dataout,
	fifo_wr_data_5,
	l1_w22_n0_mux_dataout,
	fifo_wr_data_6,
	l1_w23_n0_mux_dataout,
	fifo_wr_data_7,
	Equal3,
	length_write1,
	control_8)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a32;
input 	ram_block1a0;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a38;
input 	ram_block1a6;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a40;
input 	ram_block1a8;
input 	ram_block1a41;
input 	ram_block1a9;
input 	ram_block1a42;
input 	ram_block1a10;
input 	ram_block1a43;
input 	ram_block1a11;
input 	ram_block1a44;
input 	ram_block1a12;
input 	ram_block1a45;
input 	ram_block1a13;
input 	ram_block1a46;
input 	ram_block1a14;
input 	ram_block1a47;
input 	ram_block1a15;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	clk;
input 	readaddress_0;
input 	readaddress_1;
input 	control_2;
input 	control_0;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	src0_valid;
input 	reset_n;
input 	in_data_reg_59;
input 	mem;
input 	in_data_reg_3;
input 	address_reg_a_0;
input 	l1_w16_n0_mux_dataout;
output 	fifo_wr_data_0;
input 	p1_control;
input 	l1_w17_n0_mux_dataout;
output 	fifo_wr_data_1;
input 	l1_w18_n0_mux_dataout;
output 	fifo_wr_data_2;
input 	l1_w19_n0_mux_dataout;
output 	fifo_wr_data_3;
input 	l1_w20_n0_mux_dataout;
output 	fifo_wr_data_4;
input 	l1_w21_n0_mux_dataout;
output 	fifo_wr_data_5;
input 	l1_w22_n0_mux_dataout;
output 	fifo_wr_data_6;
input 	l1_w23_n0_mux_dataout;
output 	fifo_wr_data_7;
input 	Equal3;
output 	length_write1;
input 	control_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~0_combout ;
wire \read_data_mux_input[0]~0_combout ;
wire \readdata_mux_select[1]~0_combout ;
wire \readdata_mux_select[0]~q ;
wire \Add0~1_combout ;
wire \read_data_mux_input[1]~1_combout ;
wire \readdata_mux_select[1]~q ;
wire \fifo_wr_data~0_combout ;
wire \Equal4~0_combout ;
wire \fifo_wr_data~1_combout ;
wire \fifo_wr_data[0]~2_combout ;
wire \fifo_wr_data[0]~3_combout ;
wire \fifo_wr_data~5_combout ;
wire \fifo_wr_data~6_combout ;
wire \fifo_wr_data[1]~7_combout ;
wire \fifo_wr_data~9_combout ;
wire \fifo_wr_data~10_combout ;
wire \fifo_wr_data[2]~11_combout ;
wire \fifo_wr_data~13_combout ;
wire \fifo_wr_data~14_combout ;
wire \fifo_wr_data[3]~15_combout ;
wire \fifo_wr_data~17_combout ;
wire \fifo_wr_data~18_combout ;
wire \fifo_wr_data[4]~19_combout ;
wire \fifo_wr_data~21_combout ;
wire \fifo_wr_data~22_combout ;
wire \fifo_wr_data[5]~23_combout ;
wire \fifo_wr_data~25_combout ;
wire \fifo_wr_data~26_combout ;
wire \fifo_wr_data[6]~27_combout ;
wire \fifo_wr_data~29_combout ;
wire \fifo_wr_data~30_combout ;
wire \fifo_wr_data[7]~31_combout ;


cyclonev_lcell_comb \fifo_wr_data[0]~4 (
	.dataa(!\fifo_wr_data~0_combout ),
	.datab(!\Equal4~0_combout ),
	.datac(!l1_w16_n0_mux_dataout),
	.datad(!\fifo_wr_data~1_combout ),
	.datae(!\fifo_wr_data[0]~2_combout ),
	.dataf(!\fifo_wr_data[0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[0]~4 .extended_lut = "off";
defparam \fifo_wr_data[0]~4 .lut_mask = 64'h57FF57FFFFFF57FF;
defparam \fifo_wr_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[1]~8 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~5_combout ),
	.datad(!l1_w17_n0_mux_dataout),
	.datae(!\fifo_wr_data~6_combout ),
	.dataf(!\fifo_wr_data[1]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[1]~8 .extended_lut = "off";
defparam \fifo_wr_data[1]~8 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[1]~8 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[2]~12 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~9_combout ),
	.datad(!l1_w18_n0_mux_dataout),
	.datae(!\fifo_wr_data~10_combout ),
	.dataf(!\fifo_wr_data[2]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[2]~12 .extended_lut = "off";
defparam \fifo_wr_data[2]~12 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[2]~12 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[3]~16 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~13_combout ),
	.datad(!l1_w19_n0_mux_dataout),
	.datae(!\fifo_wr_data~14_combout ),
	.dataf(!\fifo_wr_data[3]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[3]~16 .extended_lut = "off";
defparam \fifo_wr_data[3]~16 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[3]~16 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[4]~20 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~17_combout ),
	.datad(!l1_w20_n0_mux_dataout),
	.datae(!\fifo_wr_data~18_combout ),
	.dataf(!\fifo_wr_data[4]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[4]~20 .extended_lut = "off";
defparam \fifo_wr_data[4]~20 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[4]~20 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[5]~24 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~21_combout ),
	.datad(!l1_w21_n0_mux_dataout),
	.datae(!\fifo_wr_data~22_combout ),
	.dataf(!\fifo_wr_data[5]~23_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[5]~24 .extended_lut = "off";
defparam \fifo_wr_data[5]~24 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[5]~24 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[6]~28 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~25_combout ),
	.datad(!l1_w22_n0_mux_dataout),
	.datae(!\fifo_wr_data~26_combout ),
	.dataf(!\fifo_wr_data[6]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[6]~28 .extended_lut = "off";
defparam \fifo_wr_data[6]~28 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[6]~28 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[7]~32 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\fifo_wr_data[0]~2_combout ),
	.datac(!\fifo_wr_data~29_combout ),
	.datad(!l1_w23_n0_mux_dataout),
	.datae(!\fifo_wr_data~30_combout ),
	.dataf(!\fifo_wr_data[7]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(fifo_wr_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[7]~32 .extended_lut = "off";
defparam \fifo_wr_data[7]~32 .lut_mask = 64'h0F5FFFFFCFDFFFFF;
defparam \fifo_wr_data[7]~32 .shared_arith = "off";

cyclonev_lcell_comb length_write(
	.dataa(!WideOr0),
	.datab(!wait_latency_counter_1),
	.datac(!in_data_reg_59),
	.datad(!mem),
	.datae(!Equal3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(length_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam length_write.extended_lut = "off";
defparam length_write.lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam length_write.shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!control_0),
	.datab(!\readdata_mux_select[0]~q ),
	.datac(!control_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6363636363636363;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \read_data_mux_input[0]~0 (
	.dataa(!in_data_reg_3),
	.datab(!p1_control),
	.datac(!readaddress_0),
	.datad(!length_write1),
	.datae(!\Add0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_data_mux_input[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_data_mux_input[0]~0 .extended_lut = "off";
defparam \read_data_mux_input[0]~0 .lut_mask = 64'h0F010FEF0F010FEF;
defparam \read_data_mux_input[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \readdata_mux_select[1]~0 (
	.dataa(!src0_valid),
	.datab(!in_data_reg_3),
	.datac(!p1_control),
	.datad(!length_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata_mux_select[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata_mux_select[1]~0 .extended_lut = "off";
defparam \readdata_mux_select[1]~0 .lut_mask = 64'hFF57FF57FF57FF57;
defparam \readdata_mux_select[1]~0 .shared_arith = "off";

dffeas \readdata_mux_select[0] (
	.clk(clk),
	.d(\read_data_mux_input[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_mux_select[1]~0_combout ),
	.q(\readdata_mux_select[0]~q ),
	.prn(vcc));
defparam \readdata_mux_select[0] .is_wysiwyg = "true";
defparam \readdata_mux_select[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!control_0),
	.datab(!\readdata_mux_select[0]~q ),
	.datac(!\readdata_mux_select[1]~q ),
	.datad(!control_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h1E0F1E0F1E0F1E0F;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \read_data_mux_input[1]~1 (
	.dataa(!in_data_reg_3),
	.datab(!p1_control),
	.datac(!readaddress_1),
	.datad(!length_write1),
	.datae(!\Add0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_data_mux_input[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_data_mux_input[1]~1 .extended_lut = "off";
defparam \read_data_mux_input[1]~1 .lut_mask = 64'h0F010FEF0F010FEF;
defparam \read_data_mux_input[1]~1 .shared_arith = "off";

dffeas \readdata_mux_select[1] (
	.clk(clk),
	.d(\read_data_mux_input[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\readdata_mux_select[1]~0_combout ),
	.q(\readdata_mux_select[1]~q ),
	.prn(vcc));
defparam \readdata_mux_select[1] .is_wysiwyg = "true";
defparam \readdata_mux_select[1] .power_up = "low";

cyclonev_lcell_comb \fifo_wr_data~0 (
	.dataa(!ram_block1a40),
	.datab(!ram_block1a8),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~0 .extended_lut = "off";
defparam \fifo_wr_data~0 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!control_0),
	.datab(!\readdata_mux_select[0]~q ),
	.datac(!\readdata_mux_select[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h0404040404040404;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~1 (
	.dataa(!ram_block1a56),
	.datab(!ram_block1a24),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~1 .extended_lut = "off";
defparam \fifo_wr_data~1 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~1 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[0]~2 (
	.dataa(!control_2),
	.datab(!control_0),
	.datac(!\readdata_mux_select[0]~q ),
	.datad(!\readdata_mux_select[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[0]~2 .extended_lut = "off";
defparam \fifo_wr_data[0]~2 .lut_mask = 64'h4555455545554555;
defparam \fifo_wr_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[0]~3 (
	.dataa(!ram_block1a32),
	.datab(!ram_block1a0),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[0]~3 .extended_lut = "off";
defparam \fifo_wr_data[0]~3 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~5 (
	.dataa(!ram_block1a41),
	.datab(!ram_block1a9),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~5 .extended_lut = "off";
defparam \fifo_wr_data~5 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~5 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~6 (
	.dataa(!ram_block1a57),
	.datab(!ram_block1a25),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~6 .extended_lut = "off";
defparam \fifo_wr_data~6 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~6 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[1]~7 (
	.dataa(!ram_block1a33),
	.datab(!ram_block1a1),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[1]~7 .extended_lut = "off";
defparam \fifo_wr_data[1]~7 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~9 (
	.dataa(!ram_block1a42),
	.datab(!ram_block1a10),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~9 .extended_lut = "off";
defparam \fifo_wr_data~9 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~9 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~10 (
	.dataa(!ram_block1a58),
	.datab(!ram_block1a26),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~10 .extended_lut = "off";
defparam \fifo_wr_data~10 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~10 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[2]~11 (
	.dataa(!ram_block1a34),
	.datab(!ram_block1a2),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[2]~11 .extended_lut = "off";
defparam \fifo_wr_data[2]~11 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[2]~11 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~13 (
	.dataa(!ram_block1a43),
	.datab(!ram_block1a11),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~13 .extended_lut = "off";
defparam \fifo_wr_data~13 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~13 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~14 (
	.dataa(!ram_block1a59),
	.datab(!ram_block1a27),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~14 .extended_lut = "off";
defparam \fifo_wr_data~14 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~14 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[3]~15 (
	.dataa(!ram_block1a35),
	.datab(!ram_block1a3),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[3]~15 .extended_lut = "off";
defparam \fifo_wr_data[3]~15 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[3]~15 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~17 (
	.dataa(!ram_block1a44),
	.datab(!ram_block1a12),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~17 .extended_lut = "off";
defparam \fifo_wr_data~17 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~17 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~18 (
	.dataa(!ram_block1a60),
	.datab(!ram_block1a28),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~18 .extended_lut = "off";
defparam \fifo_wr_data~18 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~18 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[4]~19 (
	.dataa(!ram_block1a36),
	.datab(!ram_block1a4),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[4]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[4]~19 .extended_lut = "off";
defparam \fifo_wr_data[4]~19 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[4]~19 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~21 (
	.dataa(!ram_block1a45),
	.datab(!ram_block1a13),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~21 .extended_lut = "off";
defparam \fifo_wr_data~21 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~21 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~22 (
	.dataa(!ram_block1a61),
	.datab(!ram_block1a29),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~22 .extended_lut = "off";
defparam \fifo_wr_data~22 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~22 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[5]~23 (
	.dataa(!ram_block1a37),
	.datab(!ram_block1a5),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[5]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[5]~23 .extended_lut = "off";
defparam \fifo_wr_data[5]~23 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[5]~23 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~25 (
	.dataa(!ram_block1a46),
	.datab(!ram_block1a14),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~25 .extended_lut = "off";
defparam \fifo_wr_data~25 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~25 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~26 (
	.dataa(!ram_block1a62),
	.datab(!ram_block1a30),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~26 .extended_lut = "off";
defparam \fifo_wr_data~26 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~26 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[6]~27 (
	.dataa(!ram_block1a38),
	.datab(!ram_block1a6),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[6]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[6]~27 .extended_lut = "off";
defparam \fifo_wr_data[6]~27 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[6]~27 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~29 (
	.dataa(!ram_block1a47),
	.datab(!ram_block1a15),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~29 .extended_lut = "off";
defparam \fifo_wr_data~29 .lut_mask = 64'h0003000000050000;
defparam \fifo_wr_data~29 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data~30 (
	.dataa(!ram_block1a63),
	.datab(!ram_block1a31),
	.datac(!control_0),
	.datad(!\readdata_mux_select[0]~q ),
	.datae(!\readdata_mux_select[1]~q ),
	.dataf(!address_reg_a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data~30 .extended_lut = "off";
defparam \fifo_wr_data~30 .lut_mask = 64'h0000000300000005;
defparam \fifo_wr_data~30 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wr_data[7]~31 (
	.dataa(!ram_block1a39),
	.datab(!ram_block1a7),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr_data[7]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr_data[7]~31 .extended_lut = "off";
defparam \fifo_wr_data[7]~31 .lut_mask = 64'h3535353535353535;
defparam \fifo_wr_data[7]~31 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	hold_waitrequest,
	WideOr0,
	wait_latency_counter_1,
	WideOr01,
	wait_latency_counter_11,
	cmd_sink_ready,
	nonposted_cmd_accepted,
	WideOr1,
	src_payload_0,
	WideOr11,
	nonposted_cmd_accepted1,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_0,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	src_data_8,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_data_13,
	src_data_14,
	src_data_15,
	src_data_16,
	src_data_17,
	src_data_18,
	src_data_19,
	src_data_20,
	src_data_21,
	src_data_22,
	src_data_23,
	src_data_24,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	src_data_29,
	src_data_30,
	src_data_31,
	src_data_881,
	src_data_891,
	src_data_901,
	src_data_911,
	src_data_921,
	src_data_931,
	src_data_941,
	src_data_951,
	src_data_961,
	src_data_971,
	src_data_981,
	src_data_991,
	altera_reset_synchronizer_int_chain_out,
	r_sync_rst,
	in_data_reg_2,
	in_data_reg_59,
	mem,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	in_data_reg_210,
	in_data_reg_591,
	mem1,
	int_nxt_addr_reg_dly_21,
	int_nxt_addr_reg_dly_41,
	int_nxt_addr_reg_dly_31,
	in_data_reg_32,
	in_data_reg_41,
	in_data_reg_51,
	in_data_reg_61,
	in_data_reg_71,
	in_data_reg_81,
	in_data_reg_91,
	in_data_reg_101,
	in_data_reg_111,
	in_data_reg_121,
	in_data_reg_131,
	in_data_reg_141,
	in_data_reg_151,
	in_data_reg_161,
	in_data_reg_171,
	in_data_reg_181,
	in_data_reg_191,
	in_data_reg_201,
	in_data_reg_211,
	in_data_reg_221,
	in_data_reg_231,
	in_data_reg_241,
	in_data_reg_251,
	in_data_reg_261,
	in_data_reg_271,
	in_data_reg_281,
	in_data_reg_291,
	in_data_reg_301,
	in_data_reg_311,
	in_data_reg_0,
	in_data_reg_1,
	dma_ctl_readdata_0,
	dma_ctl_readdata_01,
	dma_ctl_readdata_1,
	dma_ctl_readdata_11,
	dma_ctl_readdata_2,
	dma_ctl_readdata_21,
	dma_ctl_readdata_3,
	dma_ctl_readdata_31,
	dma_ctl_readdata_4,
	dma_ctl_readdata_41,
	dma_ctl_readdata_5,
	dma_ctl_readdata_51,
	dma_ctl_readdata_6,
	dma_ctl_readdata_61,
	dma_ctl_readdata_7,
	dma_ctl_readdata_71,
	dma_ctl_readdata_8,
	dma_ctl_readdata_81,
	dma_ctl_readdata_9,
	dma_ctl_readdata_91,
	dma_ctl_readdata_10,
	dma_ctl_readdata_101,
	dma_ctl_readdata_111,
	dma_ctl_readdata_112,
	dma_ctl_readdata_12,
	dma_ctl_readdata_121,
	dma_ctl_readdata_13,
	dma_ctl_readdata_131,
	dma_ctl_readdata_14,
	dma_ctl_readdata_141,
	dma_ctl_readdata_15,
	dma_ctl_readdata_151,
	dma_ctl_readdata_16,
	dma_ctl_readdata_161,
	dma_ctl_readdata_17,
	dma_ctl_readdata_171,
	dma_ctl_readdata_18,
	dma_ctl_readdata_181,
	dma_ctl_readdata_19,
	dma_ctl_readdata_191,
	dma_ctl_readdata_20,
	dma_ctl_readdata_201,
	dma_ctl_readdata_211,
	dma_ctl_readdata_212,
	dma_ctl_readdata_22,
	dma_ctl_readdata_221,
	dma_ctl_readdata_23,
	dma_ctl_readdata_231,
	dma_ctl_readdata_24,
	dma_ctl_readdata_241,
	dma_ctl_readdata_25,
	dma_ctl_readdata_251,
	dma_ctl_readdata_26,
	dma_ctl_readdata_261,
	dma_ctl_readdata_27,
	dma_ctl_readdata_271,
	dma_ctl_readdata_28,
	dma_ctl_readdata_281,
	dma_ctl_readdata_29,
	dma_ctl_readdata_291,
	dma_ctl_readdata_30,
	dma_ctl_readdata_301,
	dma_ctl_readdata_311,
	dma_ctl_readdata_312,
	in_data_reg_01,
	in_data_reg_110)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARADDR_5;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	hold_waitrequest;
output 	WideOr0;
output 	wait_latency_counter_1;
output 	WideOr01;
output 	wait_latency_counter_11;
output 	cmd_sink_ready;
output 	nonposted_cmd_accepted;
output 	WideOr1;
output 	src_payload_0;
output 	WideOr11;
output 	nonposted_cmd_accepted1;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_0;
output 	src_data_1;
output 	src_data_2;
output 	src_data_3;
output 	src_data_4;
output 	src_data_5;
output 	src_data_6;
output 	src_data_7;
output 	src_data_8;
output 	src_data_9;
output 	src_data_10;
output 	src_data_11;
output 	src_data_12;
output 	src_data_13;
output 	src_data_14;
output 	src_data_15;
output 	src_data_16;
output 	src_data_17;
output 	src_data_18;
output 	src_data_19;
output 	src_data_20;
output 	src_data_21;
output 	src_data_22;
output 	src_data_23;
output 	src_data_24;
output 	src_data_25;
output 	src_data_26;
output 	src_data_27;
output 	src_data_28;
output 	src_data_29;
output 	src_data_30;
output 	src_data_31;
output 	src_data_881;
output 	src_data_891;
output 	src_data_901;
output 	src_data_911;
output 	src_data_921;
output 	src_data_931;
output 	src_data_941;
output 	src_data_951;
output 	src_data_961;
output 	src_data_971;
output 	src_data_981;
output 	src_data_991;
input 	altera_reset_synchronizer_int_chain_out;
input 	r_sync_rst;
output 	in_data_reg_2;
output 	in_data_reg_59;
output 	mem;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
output 	in_data_reg_210;
output 	in_data_reg_591;
output 	mem1;
output 	int_nxt_addr_reg_dly_21;
output 	int_nxt_addr_reg_dly_41;
output 	int_nxt_addr_reg_dly_31;
output 	in_data_reg_32;
output 	in_data_reg_41;
output 	in_data_reg_51;
output 	in_data_reg_61;
output 	in_data_reg_71;
output 	in_data_reg_81;
output 	in_data_reg_91;
output 	in_data_reg_101;
output 	in_data_reg_111;
output 	in_data_reg_121;
output 	in_data_reg_131;
output 	in_data_reg_141;
output 	in_data_reg_151;
output 	in_data_reg_161;
output 	in_data_reg_171;
output 	in_data_reg_181;
output 	in_data_reg_191;
output 	in_data_reg_201;
output 	in_data_reg_211;
output 	in_data_reg_221;
output 	in_data_reg_231;
output 	in_data_reg_241;
output 	in_data_reg_251;
output 	in_data_reg_261;
output 	in_data_reg_271;
output 	in_data_reg_281;
output 	in_data_reg_291;
output 	in_data_reg_301;
output 	in_data_reg_311;
output 	in_data_reg_0;
output 	in_data_reg_1;
input 	dma_ctl_readdata_0;
input 	dma_ctl_readdata_01;
input 	dma_ctl_readdata_1;
input 	dma_ctl_readdata_11;
input 	dma_ctl_readdata_2;
input 	dma_ctl_readdata_21;
input 	dma_ctl_readdata_3;
input 	dma_ctl_readdata_31;
input 	dma_ctl_readdata_4;
input 	dma_ctl_readdata_41;
input 	dma_ctl_readdata_5;
input 	dma_ctl_readdata_51;
input 	dma_ctl_readdata_6;
input 	dma_ctl_readdata_61;
input 	dma_ctl_readdata_7;
input 	dma_ctl_readdata_71;
input 	dma_ctl_readdata_8;
input 	dma_ctl_readdata_81;
input 	dma_ctl_readdata_9;
input 	dma_ctl_readdata_91;
input 	dma_ctl_readdata_10;
input 	dma_ctl_readdata_101;
input 	dma_ctl_readdata_111;
input 	dma_ctl_readdata_112;
input 	dma_ctl_readdata_12;
input 	dma_ctl_readdata_121;
input 	dma_ctl_readdata_13;
input 	dma_ctl_readdata_131;
input 	dma_ctl_readdata_14;
input 	dma_ctl_readdata_141;
input 	dma_ctl_readdata_15;
input 	dma_ctl_readdata_151;
input 	dma_ctl_readdata_16;
input 	dma_ctl_readdata_161;
input 	dma_ctl_readdata_17;
input 	dma_ctl_readdata_171;
input 	dma_ctl_readdata_18;
input 	dma_ctl_readdata_181;
input 	dma_ctl_readdata_19;
input 	dma_ctl_readdata_191;
input 	dma_ctl_readdata_20;
input 	dma_ctl_readdata_201;
input 	dma_ctl_readdata_211;
input 	dma_ctl_readdata_212;
input 	dma_ctl_readdata_22;
input 	dma_ctl_readdata_221;
input 	dma_ctl_readdata_23;
input 	dma_ctl_readdata_231;
input 	dma_ctl_readdata_24;
input 	dma_ctl_readdata_241;
input 	dma_ctl_readdata_25;
input 	dma_ctl_readdata_251;
input 	dma_ctl_readdata_26;
input 	dma_ctl_readdata_261;
input 	dma_ctl_readdata_27;
input 	dma_ctl_readdata_271;
input 	dma_ctl_readdata_28;
input 	dma_ctl_readdata_281;
input 	dma_ctl_readdata_29;
input 	dma_ctl_readdata_291;
input 	dma_ctl_readdata_30;
input 	dma_ctl_readdata_301;
input 	dma_ctl_readdata_311;
input 	dma_ctl_readdata_312;
output 	in_data_reg_01;
output 	in_data_reg_110;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \dma_2_control_port_slave_translator|read_latency_shift_reg~0_combout ;
wire \dma_2_control_port_slave_agent|cp_ready~0_combout ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \dma_1_control_port_slave_translator|read_latency_shift_reg~0_combout ;
wire \dma_1_control_port_slave_agent|cp_ready~0_combout ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \cmd_demux_001|WideOr0~0_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \cmd_demux_001|WideOr0~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_rd_limiter|last_dest_id[0]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ;
wire \cmd_mux_001|saved_grant[0]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ;
wire \cmd_demux|WideOr0~0_combout ;
wire \cmd_mux|saved_grant[0]~q ;
wire \cmd_demux|WideOr0~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ;
wire \dma_1_control_port_slave_translator|read_latency_shift_reg[0]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem_used[0]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][112]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem_used[0]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][59]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][57]~q ;
wire \rsp_demux|src0_valid~combout ;
wire \dma_2_control_port_slave_translator|read_latency_shift_reg[0]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem_used[0]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][112]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem_used[0]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][59]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][57]~q ;
wire \rsp_demux_001|src0_valid~combout ;
wire \rsp_demux|src1_valid~0_combout ;
wire \dma_1_control_port_slave_agent|comb~0_combout ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][113]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][65]~q ;
wire \dma_1_control_port_slave_agent|uncompressor|last_packet_beat~0_combout ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][69]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][66]~q ;
wire \dma_1_control_port_slave_agent|uncompressor|last_packet_beat~1_combout ;
wire \rsp_mux_001|src_payload~0_combout ;
wire \rsp_demux_001|src1_valid~0_combout ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][113]~q ;
wire \dma_2_control_port_slave_agent|comb~0_combout ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][69]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][66]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][65]~q ;
wire \dma_2_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][88]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][88]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][89]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][89]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][90]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][90]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][91]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][91]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][92]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][92]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][93]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][93]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][94]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][94]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][95]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][95]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][96]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][96]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][97]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][97]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][98]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][98]~q ;
wire \dma_1_control_port_slave_agent_rsp_fifo|mem[0][99]~q ;
wire \dma_2_control_port_slave_agent_rsp_fifo|mem[0][99]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[0]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][0]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[0]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][0]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[1]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][1]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[1]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][1]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[2]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][2]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[2]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][2]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[3]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][3]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[3]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][3]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[4]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][4]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[4]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][4]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[5]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][5]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[5]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][5]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[6]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][6]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[6]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][6]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[7]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][7]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[7]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][7]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[8]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][8]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[8]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][8]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[9]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][9]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[9]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][9]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[10]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][10]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[10]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][10]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[11]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][11]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[11]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][11]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[12]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][12]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[12]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][12]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[13]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][13]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[13]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][13]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[14]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][14]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[14]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][14]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[15]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][15]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[15]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][15]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[16]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][16]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[16]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][16]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[17]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][17]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[17]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][17]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[18]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][18]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[18]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][18]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[19]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][19]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[19]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][19]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[20]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][20]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[20]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][20]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[21]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][21]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[21]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][21]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[22]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][22]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[22]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][22]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[23]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][23]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[23]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][23]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[24]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][24]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[24]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][24]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[25]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][25]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[25]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][25]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[26]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][26]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[26]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][26]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[27]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][27]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[27]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][27]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[28]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][28]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[28]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][28]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[29]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][29]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[29]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][29]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[30]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][30]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[30]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][30]~q ;
wire \dma_1_control_port_slave_translator|av_readdata_pre[31]~q ;
wire \dma_1_control_port_slave_agent_rdata_fifo|mem[0][31]~q ;
wire \dma_2_control_port_slave_translator|av_readdata_pre[31]~q ;
wire \dma_2_control_port_slave_agent_rdata_fifo|mem[0][31]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~0_combout ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \dma_2_control_port_slave_agent|cp_ready~2_combout ;
wire \rsp_demux_001|WideOr0~0_combout ;
wire \dma_2_control_port_slave_agent_rsp_fifo|read~0_combout ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \cmd_mux_001|src_data[78]~combout ;
wire \cmd_mux_001|src_data[79]~combout ;
wire \cmd_mux_001|src_data[35]~combout ;
wire \cmd_mux_001|src_data[34]~combout ;
wire \cmd_mux_001|src_data[33]~combout ;
wire \cmd_mux_001|src_data[32]~combout ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~1_combout ;
wire \cmd_mux_001|src_payload[0]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~4_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add2~1_combout ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~2_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \dma_1_control_port_slave_agent|cp_ready~2_combout ;
wire \dma_1_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ;
wire \rsp_demux|WideOr0~0_combout ;
wire \dma_1_control_port_slave_agent_rsp_fifo|read~0_combout ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \cmd_mux|src_data[78]~combout ;
wire \cmd_mux|src_data[79]~combout ;
wire \cmd_mux|src_data[35]~combout ;
wire \cmd_mux|src_data[34]~combout ;
wire \cmd_mux|src_data[33]~combout ;
wire \cmd_mux|src_data[32]~combout ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~3_combout ;
wire \cmd_mux|src_payload[0]~combout ;
wire \cmd_demux_001|WideOr0~2_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[5]~0_combout ;
wire \dma_1_control_port_slave_agent|rp_valid~combout ;
wire \dma_2_control_port_slave_agent|rp_valid~combout ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \cmd_mux|src_payload~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector4~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector11~1_combout ;
wire \cmd_mux|src_data[72]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[4]~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector2~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector9~1_combout ;
wire \cmd_mux|src_data[74]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~2_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector3~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector10~1_combout ;
wire \cmd_mux|src_data[73]~combout ;
wire \cmd_mux|src_payload~1_combout ;
wire \cmd_mux|src_payload~2_combout ;
wire \cmd_mux|src_payload~3_combout ;
wire \cmd_mux|src_payload~4_combout ;
wire \cmd_mux|src_payload~5_combout ;
wire \cmd_mux|src_payload~6_combout ;
wire \cmd_mux|src_payload~7_combout ;
wire \cmd_mux|src_payload~8_combout ;
wire \cmd_mux|src_payload~9_combout ;
wire \cmd_mux|src_payload~10_combout ;
wire \cmd_mux|src_payload~11_combout ;
wire \cmd_mux|src_payload~12_combout ;
wire \cmd_mux|src_payload~13_combout ;
wire \cmd_mux|src_payload~14_combout ;
wire \cmd_mux|src_payload~15_combout ;
wire \cmd_mux|src_payload~16_combout ;
wire \cmd_mux|src_payload~17_combout ;
wire \cmd_mux|src_payload~18_combout ;
wire \cmd_mux|src_payload~19_combout ;
wire \cmd_mux|src_payload~20_combout ;
wire \cmd_mux|src_payload~21_combout ;
wire \cmd_mux|src_payload~22_combout ;
wire \cmd_mux|src_payload~23_combout ;
wire \cmd_mux|src_payload~24_combout ;
wire \cmd_mux|src_payload~25_combout ;
wire \cmd_mux|src_payload~26_combout ;
wire \cmd_mux|src_payload~27_combout ;
wire \cmd_mux|src_payload~28_combout ;
wire \cmd_mux|src_payload~29_combout ;
wire \cmd_mux_001|src_payload~0_combout ;
wire \cmd_mux_001|src_data[72]~combout ;
wire \cmd_mux_001|src_data[74]~combout ;
wire \cmd_mux_001|src_data[73]~combout ;
wire \cmd_mux_001|src_payload~1_combout ;
wire \cmd_mux_001|src_payload~2_combout ;
wire \cmd_mux_001|src_payload~3_combout ;
wire \cmd_mux_001|src_payload~4_combout ;
wire \cmd_mux_001|src_payload~5_combout ;
wire \cmd_mux_001|src_payload~6_combout ;
wire \cmd_mux_001|src_payload~7_combout ;
wire \cmd_mux_001|src_payload~8_combout ;
wire \cmd_mux_001|src_payload~9_combout ;
wire \cmd_mux_001|src_payload~10_combout ;
wire \cmd_mux_001|src_payload~11_combout ;
wire \cmd_mux_001|src_payload~12_combout ;
wire \cmd_mux_001|src_payload~13_combout ;
wire \cmd_mux_001|src_payload~14_combout ;
wire \cmd_mux_001|src_payload~15_combout ;
wire \cmd_mux_001|src_payload~16_combout ;
wire \cmd_mux_001|src_payload~17_combout ;
wire \cmd_mux_001|src_payload~18_combout ;
wire \cmd_mux_001|src_payload~19_combout ;
wire \cmd_mux_001|src_payload~20_combout ;
wire \cmd_mux_001|src_payload~21_combout ;
wire \cmd_mux_001|src_payload~22_combout ;
wire \cmd_mux_001|src_payload~23_combout ;
wire \cmd_mux_001|src_payload~24_combout ;
wire \cmd_mux_001|src_payload~25_combout ;
wire \cmd_mux_001|src_payload~26_combout ;
wire \cmd_mux_001|src_payload~27_combout ;
wire \cmd_mux_001|src_payload~28_combout ;
wire \cmd_mux_001|src_payload~29_combout ;
wire \cmd_mux_001|src_payload~30_combout ;
wire \cmd_mux_001|src_payload~31_combout ;
wire \cmd_demux|WideOr0~2_combout ;
wire \cmd_demux|WideOr0~3_combout ;
wire \cmd_mux|src_data[88]~combout ;
wire \cmd_mux_001|src_data[88]~combout ;
wire \cmd_mux|src_data[89]~combout ;
wire \cmd_mux_001|src_data[89]~combout ;
wire \cmd_mux|src_data[90]~combout ;
wire \cmd_mux_001|src_data[90]~combout ;
wire \cmd_mux|src_data[91]~combout ;
wire \cmd_mux_001|src_data[91]~combout ;
wire \cmd_mux|src_data[92]~combout ;
wire \cmd_mux_001|src_data[92]~combout ;
wire \cmd_mux|src_data[93]~combout ;
wire \cmd_mux_001|src_data[93]~combout ;
wire \cmd_mux|src_data[94]~combout ;
wire \cmd_mux_001|src_data[94]~combout ;
wire \cmd_mux|src_data[95]~combout ;
wire \cmd_mux_001|src_data[95]~combout ;
wire \cmd_mux|src_data[96]~combout ;
wire \cmd_mux_001|src_data[96]~combout ;
wire \cmd_mux|src_data[97]~combout ;
wire \cmd_mux_001|src_data[97]~combout ;
wire \cmd_mux|src_data[98]~combout ;
wire \cmd_mux_001|src_data[98]~combout ;
wire \cmd_mux|src_data[99]~combout ;
wire \cmd_mux_001|src_data[99]~combout ;
wire \cmd_mux|src_payload~30_combout ;
wire \cmd_mux|src_payload~31_combout ;
wire \cmd_mux|src_data[77]~combout ;
wire \cmd_mux_001|src_data[77]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector5~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector12~1_combout ;
wire \cmd_mux|src_data[71]~combout ;
wire \cmd_mux_001|src_data[71]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~2_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector6~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Selector13~1_combout ;
wire \cmd_mux|src_data[70]~combout ;
wire \cmd_mux_001|src_data[70]~combout ;


Computer_System_altera_merlin_slave_translator_1 dma_2_control_port_slave_translator(
	.clk(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.WideOr0(WideOr0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.read_latency_shift_reg(\dma_2_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg_0(\dma_2_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\dma_2_control_port_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\dma_2_control_port_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\dma_2_control_port_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\dma_2_control_port_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\dma_2_control_port_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\dma_2_control_port_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\dma_2_control_port_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\dma_2_control_port_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\dma_2_control_port_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\dma_2_control_port_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\dma_2_control_port_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\dma_2_control_port_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\dma_2_control_port_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\dma_2_control_port_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\dma_2_control_port_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\dma_2_control_port_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\dma_2_control_port_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\dma_2_control_port_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\dma_2_control_port_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\dma_2_control_port_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_20(\dma_2_control_port_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\dma_2_control_port_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\dma_2_control_port_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\dma_2_control_port_slave_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\dma_2_control_port_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\dma_2_control_port_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\dma_2_control_port_slave_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\dma_2_control_port_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\dma_2_control_port_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\dma_2_control_port_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\dma_2_control_port_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\dma_2_control_port_slave_translator|av_readdata_pre[31]~q ),
	.reset(r_sync_rst),
	.in_data_reg_59(in_data_reg_591),
	.mem(mem1),
	.in_data_reg_60(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.av_readdata({dma_ctl_readdata_312,dma_ctl_readdata_301,dma_ctl_readdata_291,dma_ctl_readdata_281,dma_ctl_readdata_271,dma_ctl_readdata_261,dma_ctl_readdata_251,dma_ctl_readdata_241,dma_ctl_readdata_231,dma_ctl_readdata_221,dma_ctl_readdata_212,dma_ctl_readdata_201,
dma_ctl_readdata_191,dma_ctl_readdata_181,dma_ctl_readdata_171,dma_ctl_readdata_161,dma_ctl_readdata_151,dma_ctl_readdata_141,dma_ctl_readdata_131,dma_ctl_readdata_121,dma_ctl_readdata_112,dma_ctl_readdata_101,dma_ctl_readdata_91,dma_ctl_readdata_81,
dma_ctl_readdata_71,dma_ctl_readdata_61,dma_ctl_readdata_51,dma_ctl_readdata_41,dma_ctl_readdata_31,dma_ctl_readdata_21,dma_ctl_readdata_11,dma_ctl_readdata_01}));

Computer_System_altera_merlin_slave_translator dma_1_control_port_slave_translator(
	.clk(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.WideOr0(WideOr01),
	.wait_latency_counter_1(wait_latency_counter_11),
	.read_latency_shift_reg(\dma_1_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg_0(\dma_1_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\dma_1_control_port_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\dma_1_control_port_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\dma_1_control_port_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\dma_1_control_port_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\dma_1_control_port_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\dma_1_control_port_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\dma_1_control_port_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\dma_1_control_port_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\dma_1_control_port_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\dma_1_control_port_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\dma_1_control_port_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\dma_1_control_port_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\dma_1_control_port_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\dma_1_control_port_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\dma_1_control_port_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\dma_1_control_port_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\dma_1_control_port_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\dma_1_control_port_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\dma_1_control_port_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\dma_1_control_port_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_20(\dma_1_control_port_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\dma_1_control_port_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\dma_1_control_port_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\dma_1_control_port_slave_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\dma_1_control_port_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\dma_1_control_port_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\dma_1_control_port_slave_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\dma_1_control_port_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\dma_1_control_port_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\dma_1_control_port_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\dma_1_control_port_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\dma_1_control_port_slave_translator|av_readdata_pre[31]~q ),
	.reset(r_sync_rst),
	.in_data_reg_59(in_data_reg_59),
	.mem(mem),
	.in_data_reg_60(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.av_readdata({dma_ctl_readdata_311,dma_ctl_readdata_30,dma_ctl_readdata_29,dma_ctl_readdata_28,dma_ctl_readdata_27,dma_ctl_readdata_26,dma_ctl_readdata_25,dma_ctl_readdata_24,dma_ctl_readdata_23,dma_ctl_readdata_22,dma_ctl_readdata_211,dma_ctl_readdata_20,dma_ctl_readdata_19,
dma_ctl_readdata_18,dma_ctl_readdata_17,dma_ctl_readdata_16,dma_ctl_readdata_15,dma_ctl_readdata_14,dma_ctl_readdata_13,dma_ctl_readdata_12,dma_ctl_readdata_111,dma_ctl_readdata_10,dma_ctl_readdata_9,dma_ctl_readdata_8,dma_ctl_readdata_7,dma_ctl_readdata_6,
dma_ctl_readdata_5,dma_ctl_readdata_4,dma_ctl_readdata_3,dma_ctl_readdata_2,dma_ctl_readdata_1,dma_ctl_readdata_0}));

Computer_System_Computer_System_mm_interconnect_0_rsp_mux_1 rsp_mux_001(
	.read_latency_shift_reg_0(\dma_1_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_1_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_57_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.read_latency_shift_reg_01(\dma_2_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_01(\dma_2_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.src1_valid(\rsp_demux|src1_valid~0_combout ),
	.comb(\dma_1_control_port_slave_agent|comb~0_combout ),
	.mem_113_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][113]~q ),
	.mem_65_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\dma_1_control_port_slave_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\dma_1_control_port_slave_agent|uncompressor|last_packet_beat~1_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.src1_valid1(\rsp_demux_001|src1_valid~0_combout ),
	.mem_113_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][113]~q ),
	.last_packet_beat2(\dma_2_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.src_payload_0(src_payload_0),
	.WideOr11(WideOr11),
	.mem_88_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][88]~q ),
	.mem_88_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][89]~q ),
	.mem_89_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][90]~q ),
	.mem_90_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][91]~q ),
	.mem_91_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][99]~q ),
	.av_readdata_pre_0(\dma_1_control_port_slave_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_01(\dma_2_control_port_slave_translator|av_readdata_pre[0]~q ),
	.mem_0_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_1(\dma_1_control_port_slave_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_11(\dma_2_control_port_slave_translator|av_readdata_pre[1]~q ),
	.mem_1_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_2(\dma_1_control_port_slave_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_21(\dma_2_control_port_slave_translator|av_readdata_pre[2]~q ),
	.mem_2_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_3(\dma_1_control_port_slave_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_31(\dma_2_control_port_slave_translator|av_readdata_pre[3]~q ),
	.mem_3_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_4(\dma_1_control_port_slave_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_41(\dma_2_control_port_slave_translator|av_readdata_pre[4]~q ),
	.mem_4_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_5(\dma_1_control_port_slave_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_51(\dma_2_control_port_slave_translator|av_readdata_pre[5]~q ),
	.mem_5_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_6(\dma_1_control_port_slave_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_61(\dma_2_control_port_slave_translator|av_readdata_pre[6]~q ),
	.mem_6_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_7(\dma_1_control_port_slave_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_71(\dma_2_control_port_slave_translator|av_readdata_pre[7]~q ),
	.mem_7_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_8(\dma_1_control_port_slave_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_81(\dma_2_control_port_slave_translator|av_readdata_pre[8]~q ),
	.mem_8_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_9(\dma_1_control_port_slave_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_91(\dma_2_control_port_slave_translator|av_readdata_pre[9]~q ),
	.mem_9_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_10(\dma_1_control_port_slave_translator|av_readdata_pre[10]~q ),
	.mem_10_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_101(\dma_2_control_port_slave_translator|av_readdata_pre[10]~q ),
	.mem_10_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][10]~q ),
	.src_data_10(src_data_10),
	.av_readdata_pre_111(\dma_1_control_port_slave_translator|av_readdata_pre[11]~q ),
	.mem_11_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_112(\dma_2_control_port_slave_translator|av_readdata_pre[11]~q ),
	.mem_11_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][11]~q ),
	.src_data_11(src_data_11),
	.av_readdata_pre_12(\dma_1_control_port_slave_translator|av_readdata_pre[12]~q ),
	.mem_12_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_121(\dma_2_control_port_slave_translator|av_readdata_pre[12]~q ),
	.mem_12_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][12]~q ),
	.src_data_12(src_data_12),
	.av_readdata_pre_13(\dma_1_control_port_slave_translator|av_readdata_pre[13]~q ),
	.mem_13_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_131(\dma_2_control_port_slave_translator|av_readdata_pre[13]~q ),
	.mem_13_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][13]~q ),
	.src_data_13(src_data_13),
	.av_readdata_pre_14(\dma_1_control_port_slave_translator|av_readdata_pre[14]~q ),
	.mem_14_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_141(\dma_2_control_port_slave_translator|av_readdata_pre[14]~q ),
	.mem_14_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_15(\dma_1_control_port_slave_translator|av_readdata_pre[15]~q ),
	.mem_15_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_151(\dma_2_control_port_slave_translator|av_readdata_pre[15]~q ),
	.mem_15_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][15]~q ),
	.src_data_15(src_data_15),
	.av_readdata_pre_16(\dma_1_control_port_slave_translator|av_readdata_pre[16]~q ),
	.mem_16_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_161(\dma_2_control_port_slave_translator|av_readdata_pre[16]~q ),
	.mem_16_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][16]~q ),
	.src_data_16(src_data_16),
	.av_readdata_pre_17(\dma_1_control_port_slave_translator|av_readdata_pre[17]~q ),
	.mem_17_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_171(\dma_2_control_port_slave_translator|av_readdata_pre[17]~q ),
	.mem_17_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][17]~q ),
	.src_data_17(src_data_17),
	.av_readdata_pre_18(\dma_1_control_port_slave_translator|av_readdata_pre[18]~q ),
	.mem_18_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_181(\dma_2_control_port_slave_translator|av_readdata_pre[18]~q ),
	.mem_18_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][18]~q ),
	.src_data_18(src_data_18),
	.av_readdata_pre_19(\dma_1_control_port_slave_translator|av_readdata_pre[19]~q ),
	.mem_19_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_191(\dma_2_control_port_slave_translator|av_readdata_pre[19]~q ),
	.mem_19_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][19]~q ),
	.src_data_19(src_data_19),
	.av_readdata_pre_20(\dma_1_control_port_slave_translator|av_readdata_pre[20]~q ),
	.mem_20_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_201(\dma_2_control_port_slave_translator|av_readdata_pre[20]~q ),
	.mem_20_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][20]~q ),
	.src_data_20(src_data_20),
	.av_readdata_pre_211(\dma_1_control_port_slave_translator|av_readdata_pre[21]~q ),
	.mem_21_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_212(\dma_2_control_port_slave_translator|av_readdata_pre[21]~q ),
	.mem_21_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][21]~q ),
	.src_data_21(src_data_21),
	.av_readdata_pre_22(\dma_1_control_port_slave_translator|av_readdata_pre[22]~q ),
	.mem_22_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_221(\dma_2_control_port_slave_translator|av_readdata_pre[22]~q ),
	.mem_22_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][22]~q ),
	.src_data_22(src_data_22),
	.av_readdata_pre_23(\dma_1_control_port_slave_translator|av_readdata_pre[23]~q ),
	.mem_23_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_231(\dma_2_control_port_slave_translator|av_readdata_pre[23]~q ),
	.mem_23_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][23]~q ),
	.src_data_23(src_data_23),
	.av_readdata_pre_24(\dma_1_control_port_slave_translator|av_readdata_pre[24]~q ),
	.mem_24_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_241(\dma_2_control_port_slave_translator|av_readdata_pre[24]~q ),
	.mem_24_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][24]~q ),
	.src_data_24(src_data_24),
	.av_readdata_pre_25(\dma_1_control_port_slave_translator|av_readdata_pre[25]~q ),
	.mem_25_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_251(\dma_2_control_port_slave_translator|av_readdata_pre[25]~q ),
	.mem_25_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][25]~q ),
	.src_data_25(src_data_25),
	.av_readdata_pre_26(\dma_1_control_port_slave_translator|av_readdata_pre[26]~q ),
	.mem_26_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_261(\dma_2_control_port_slave_translator|av_readdata_pre[26]~q ),
	.mem_26_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][26]~q ),
	.src_data_26(src_data_26),
	.av_readdata_pre_27(\dma_1_control_port_slave_translator|av_readdata_pre[27]~q ),
	.mem_27_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_271(\dma_2_control_port_slave_translator|av_readdata_pre[27]~q ),
	.mem_27_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][27]~q ),
	.src_data_27(src_data_27),
	.av_readdata_pre_28(\dma_1_control_port_slave_translator|av_readdata_pre[28]~q ),
	.mem_28_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_281(\dma_2_control_port_slave_translator|av_readdata_pre[28]~q ),
	.mem_28_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][28]~q ),
	.src_data_28(src_data_28),
	.av_readdata_pre_29(\dma_1_control_port_slave_translator|av_readdata_pre[29]~q ),
	.mem_29_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_291(\dma_2_control_port_slave_translator|av_readdata_pre[29]~q ),
	.mem_29_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][29]~q ),
	.src_data_29(src_data_29),
	.av_readdata_pre_30(\dma_1_control_port_slave_translator|av_readdata_pre[30]~q ),
	.mem_30_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_301(\dma_2_control_port_slave_translator|av_readdata_pre[30]~q ),
	.mem_30_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][30]~q ),
	.src_data_30(src_data_30),
	.av_readdata_pre_311(\dma_1_control_port_slave_translator|av_readdata_pre[31]~q ),
	.mem_31_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][31]~q ),
	.av_readdata_pre_312(\dma_2_control_port_slave_translator|av_readdata_pre[31]~q ),
	.mem_31_01(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][31]~q ),
	.src_data_31(src_data_31),
	.src_data_88(src_data_881),
	.src_data_89(src_data_891),
	.src_data_90(src_data_901),
	.src_data_91(src_data_911),
	.src_data_92(src_data_921),
	.src_data_93(src_data_931),
	.src_data_94(src_data_941),
	.src_data_95(src_data_951),
	.src_data_96(src_data_961),
	.src_data_97(src_data_971),
	.src_data_98(src_data_981),
	.src_data_99(src_data_991));

Computer_System_Computer_System_mm_interconnect_0_rsp_mux rsp_mux(
	.src0_valid(\rsp_demux|src0_valid~combout ),
	.src0_valid1(\rsp_demux_001|src0_valid~combout ),
	.WideOr11(WideOr1),
	.mem_88_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][88]~q ),
	.mem_88_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][88]~q ),
	.src_data_88(src_data_88),
	.mem_89_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][89]~q ),
	.mem_89_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][89]~q ),
	.src_data_89(src_data_89),
	.mem_90_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][90]~q ),
	.mem_90_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][90]~q ),
	.src_data_90(src_data_90),
	.mem_91_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][91]~q ),
	.mem_91_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][91]~q ),
	.src_data_91(src_data_91),
	.mem_92_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][92]~q ),
	.src_data_92(src_data_92),
	.mem_93_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][93]~q ),
	.src_data_93(src_data_93),
	.mem_94_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][94]~q ),
	.src_data_94(src_data_94),
	.mem_95_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][95]~q ),
	.src_data_95(src_data_95),
	.mem_96_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][96]~q ),
	.src_data_96(src_data_96),
	.mem_97_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][97]~q ),
	.src_data_97(src_data_97),
	.mem_98_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][98]~q ),
	.src_data_98(src_data_98),
	.mem_99_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_01(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][99]~q ),
	.src_data_99(src_data_99));

Computer_System_Computer_System_mm_interconnect_0_rsp_demux_1 rsp_demux_001(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\dma_2_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_2_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux_001|src0_valid~combout ),
	.src1_valid(\rsp_demux_001|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_001|WideOr0~0_combout ));

Computer_System_Computer_System_mm_interconnect_0_rsp_demux rsp_demux(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\dma_1_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_1_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux|src0_valid~combout ),
	.src1_valid(\rsp_demux|src1_valid~0_combout ),
	.WideOr0(\rsp_demux|WideOr0~0_combout ));

Computer_System_Computer_System_mm_interconnect_0_cmd_mux_1 cmd_mux_001(
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.outclk_wire_0(outclk_wire_0),
	.nxt_in_ready(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.awready(\arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.r_sync_rst(r_sync_rst),
	.cmd_src_valid_1(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.src_data_78(\cmd_mux_001|src_data[78]~combout ),
	.src_data_79(\cmd_mux_001|src_data[79]~combout ),
	.src_data_35(\cmd_mux_001|src_data[35]~combout ),
	.src_data_34(\cmd_mux_001|src_data[34]~combout ),
	.src_data_33(\cmd_mux_001|src_data[33]~combout ),
	.src_data_32(\cmd_mux_001|src_data[32]~combout ),
	.cmd_src_valid_11(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~1_combout ),
	.src_payload_0(\cmd_mux_001|src_payload[0]~combout ),
	.Selector4(\arm_a9_hps_h2f_lw_axi_master_agent|Selector4~0_combout ),
	.Selector11(\arm_a9_hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.Selector2(\arm_a9_hps_h2f_lw_axi_master_agent|Selector2~0_combout ),
	.Selector9(\arm_a9_hps_h2f_lw_axi_master_agent|Selector9~1_combout ),
	.Selector3(\arm_a9_hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\arm_a9_hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_data_72(\cmd_mux_001|src_data[72]~combout ),
	.src_data_74(\cmd_mux_001|src_data[74]~combout ),
	.src_data_73(\cmd_mux_001|src_data[73]~combout ),
	.src_payload1(\cmd_mux_001|src_payload~1_combout ),
	.src_payload2(\cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\cmd_mux_001|src_payload~3_combout ),
	.src_payload4(\cmd_mux_001|src_payload~4_combout ),
	.src_payload5(\cmd_mux_001|src_payload~5_combout ),
	.src_payload6(\cmd_mux_001|src_payload~6_combout ),
	.src_payload7(\cmd_mux_001|src_payload~7_combout ),
	.src_payload8(\cmd_mux_001|src_payload~8_combout ),
	.src_payload9(\cmd_mux_001|src_payload~9_combout ),
	.src_payload10(\cmd_mux_001|src_payload~10_combout ),
	.src_payload11(\cmd_mux_001|src_payload~11_combout ),
	.src_payload12(\cmd_mux_001|src_payload~12_combout ),
	.src_payload13(\cmd_mux_001|src_payload~13_combout ),
	.src_payload14(\cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\cmd_mux_001|src_payload~15_combout ),
	.src_payload16(\cmd_mux_001|src_payload~16_combout ),
	.src_payload17(\cmd_mux_001|src_payload~17_combout ),
	.src_payload18(\cmd_mux_001|src_payload~18_combout ),
	.src_payload19(\cmd_mux_001|src_payload~19_combout ),
	.src_payload20(\cmd_mux_001|src_payload~20_combout ),
	.src_payload21(\cmd_mux_001|src_payload~21_combout ),
	.src_payload22(\cmd_mux_001|src_payload~22_combout ),
	.src_payload23(\cmd_mux_001|src_payload~23_combout ),
	.src_payload24(\cmd_mux_001|src_payload~24_combout ),
	.src_payload25(\cmd_mux_001|src_payload~25_combout ),
	.src_payload26(\cmd_mux_001|src_payload~26_combout ),
	.src_payload27(\cmd_mux_001|src_payload~27_combout ),
	.src_payload28(\cmd_mux_001|src_payload~28_combout ),
	.src_payload29(\cmd_mux_001|src_payload~29_combout ),
	.src_payload30(\cmd_mux_001|src_payload~30_combout ),
	.src_payload31(\cmd_mux_001|src_payload~31_combout ),
	.src_data_88(\cmd_mux_001|src_data[88]~combout ),
	.src_data_89(\cmd_mux_001|src_data[89]~combout ),
	.src_data_90(\cmd_mux_001|src_data[90]~combout ),
	.src_data_91(\cmd_mux_001|src_data[91]~combout ),
	.src_data_92(\cmd_mux_001|src_data[92]~combout ),
	.src_data_93(\cmd_mux_001|src_data[93]~combout ),
	.src_data_94(\cmd_mux_001|src_data[94]~combout ),
	.src_data_95(\cmd_mux_001|src_data[95]~combout ),
	.src_data_96(\cmd_mux_001|src_data[96]~combout ),
	.src_data_97(\cmd_mux_001|src_data[97]~combout ),
	.src_data_98(\cmd_mux_001|src_data[98]~combout ),
	.src_data_99(\cmd_mux_001|src_data[99]~combout ),
	.src_data_77(\cmd_mux_001|src_data[77]~combout ),
	.Selector5(\arm_a9_hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Selector12(\arm_a9_hps_h2f_lw_axi_master_agent|Selector12~1_combout ),
	.src_data_71(\cmd_mux_001|src_data[71]~combout ),
	.Selector6(\arm_a9_hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.Selector13(\arm_a9_hps_h2f_lw_axi_master_agent|Selector13~1_combout ),
	.src_data_70(\cmd_mux_001|src_data[70]~combout ));

Computer_System_Computer_System_mm_interconnect_0_cmd_mux cmd_mux(
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.outclk_wire_0(outclk_wire_0),
	.nxt_in_ready(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.awready(\arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.r_sync_rst(r_sync_rst),
	.cmd_src_valid_0(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~2_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.cmd_src_valid_01(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~3_combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.Selector4(\arm_a9_hps_h2f_lw_axi_master_agent|Selector4~0_combout ),
	.Selector11(\arm_a9_hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.src_data_72(\cmd_mux|src_data[72]~combout ),
	.Selector2(\arm_a9_hps_h2f_lw_axi_master_agent|Selector2~0_combout ),
	.Selector9(\arm_a9_hps_h2f_lw_axi_master_agent|Selector9~1_combout ),
	.src_data_74(\cmd_mux|src_data[74]~combout ),
	.Selector3(\arm_a9_hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\arm_a9_hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.src_data_73(\cmd_mux|src_data[73]~combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.src_payload3(\cmd_mux|src_payload~3_combout ),
	.src_payload4(\cmd_mux|src_payload~4_combout ),
	.src_payload5(\cmd_mux|src_payload~5_combout ),
	.src_payload6(\cmd_mux|src_payload~6_combout ),
	.src_payload7(\cmd_mux|src_payload~7_combout ),
	.src_payload8(\cmd_mux|src_payload~8_combout ),
	.src_payload9(\cmd_mux|src_payload~9_combout ),
	.src_payload10(\cmd_mux|src_payload~10_combout ),
	.src_payload11(\cmd_mux|src_payload~11_combout ),
	.src_payload12(\cmd_mux|src_payload~12_combout ),
	.src_payload13(\cmd_mux|src_payload~13_combout ),
	.src_payload14(\cmd_mux|src_payload~14_combout ),
	.src_payload15(\cmd_mux|src_payload~15_combout ),
	.src_payload16(\cmd_mux|src_payload~16_combout ),
	.src_payload17(\cmd_mux|src_payload~17_combout ),
	.src_payload18(\cmd_mux|src_payload~18_combout ),
	.src_payload19(\cmd_mux|src_payload~19_combout ),
	.src_payload20(\cmd_mux|src_payload~20_combout ),
	.src_payload21(\cmd_mux|src_payload~21_combout ),
	.src_payload22(\cmd_mux|src_payload~22_combout ),
	.src_payload23(\cmd_mux|src_payload~23_combout ),
	.src_payload24(\cmd_mux|src_payload~24_combout ),
	.src_payload25(\cmd_mux|src_payload~25_combout ),
	.src_payload26(\cmd_mux|src_payload~26_combout ),
	.src_payload27(\cmd_mux|src_payload~27_combout ),
	.src_payload28(\cmd_mux|src_payload~28_combout ),
	.src_payload29(\cmd_mux|src_payload~29_combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.src_payload30(\cmd_mux|src_payload~30_combout ),
	.src_payload31(\cmd_mux|src_payload~31_combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.Selector5(\arm_a9_hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Selector12(\arm_a9_hps_h2f_lw_axi_master_agent|Selector12~1_combout ),
	.src_data_71(\cmd_mux|src_data[71]~combout ),
	.Selector6(\arm_a9_hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.Selector13(\arm_a9_hps_h2f_lw_axi_master_agent|Selector13~1_combout ),
	.src_data_70(\cmd_mux|src_data[70]~combout ));

Computer_System_Computer_System_mm_interconnect_0_cmd_demux_1 cmd_demux_001(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARADDR_5(h2f_lw_ARADDR_5),
	.nxt_in_ready(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.WideOr0(\cmd_demux_001|WideOr0~0_combout ),
	.saved_grant_11(\cmd_mux|saved_grant[1]~q ),
	.WideOr01(\cmd_demux_001|WideOr0~1_combout ),
	.last_dest_id_0(\arm_a9_hps_h2f_lw_axi_master_rd_limiter|last_dest_id[0]~q ),
	.has_pending_responses(\arm_a9_hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.last_channel_0(\arm_a9_hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.WideOr02(\cmd_demux_001|WideOr0~2_combout ));

Computer_System_Computer_System_mm_interconnect_0_cmd_demux cmd_demux(
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.nxt_in_ready(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.sop_enable(\arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_5(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.saved_grant_01(\cmd_mux|saved_grant[0]~q ),
	.WideOr01(\cmd_demux|WideOr0~1_combout ),
	.WideOr02(\cmd_demux|WideOr0~2_combout ),
	.WideOr03(\cmd_demux|WideOr0~3_combout ));

Computer_System_altera_merlin_burst_adapter_1 dma_2_control_port_slave_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.outclk_wire_0(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.stateST_COMP_TRANS(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(WideOr0),
	.read_latency_shift_reg(\dma_2_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.cp_ready(\dma_2_control_port_slave_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.sop_enable(\arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.awready(\arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.r_sync_rst(r_sync_rst),
	.in_data_reg_2(in_data_reg_210),
	.in_data_reg_59(in_data_reg_591),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_21),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_41),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_31),
	.in_data_reg_3(in_data_reg_32),
	.in_data_reg_4(in_data_reg_41),
	.in_data_reg_5(in_data_reg_51),
	.in_data_reg_6(in_data_reg_61),
	.in_data_reg_7(in_data_reg_71),
	.in_data_reg_8(in_data_reg_81),
	.in_data_reg_9(in_data_reg_91),
	.in_data_reg_10(in_data_reg_101),
	.in_data_reg_11(in_data_reg_111),
	.in_data_reg_12(in_data_reg_121),
	.in_data_reg_13(in_data_reg_131),
	.in_data_reg_14(in_data_reg_141),
	.in_data_reg_15(in_data_reg_151),
	.in_data_reg_16(in_data_reg_161),
	.in_data_reg_17(in_data_reg_171),
	.in_data_reg_18(in_data_reg_181),
	.in_data_reg_19(in_data_reg_191),
	.in_data_reg_20(in_data_reg_201),
	.in_data_reg_21(in_data_reg_211),
	.in_data_reg_22(in_data_reg_221),
	.in_data_reg_23(in_data_reg_231),
	.in_data_reg_24(in_data_reg_241),
	.in_data_reg_25(in_data_reg_251),
	.in_data_reg_26(in_data_reg_261),
	.in_data_reg_27(in_data_reg_271),
	.in_data_reg_28(in_data_reg_281),
	.in_data_reg_29(in_data_reg_291),
	.in_data_reg_30(in_data_reg_301),
	.in_data_reg_31(in_data_reg_311),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.nxt_out_eop(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.cmd_src_valid_1(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.cp_ready1(\dma_2_control_port_slave_agent|cp_ready~2_combout ),
	.in_data_reg_60(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux_001|src_data[78]~combout ),
	.src_data_79(\cmd_mux_001|src_data[79]~combout ),
	.src_data_35(\cmd_mux_001|src_data[35]~combout ),
	.src_data_34(\cmd_mux_001|src_data[34]~combout ),
	.src_data_33(\cmd_mux_001|src_data[33]~combout ),
	.src_data_32(\cmd_mux_001|src_data[32]~combout ),
	.out_uncomp_byte_cnt_reg_6(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_byte_cnt_reg_2(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cmd_src_valid_11(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~1_combout ),
	.src_payload_0(\cmd_mux_001|src_payload[0]~combout ),
	.burst_bytecount_2(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~0_combout ),
	.burst_bytecount_3(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ),
	.burst_bytecount_4(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.burst_bytecount_5(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ),
	.Add2(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.burst_bytecount_6(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~4_combout ),
	.Add21(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.WideNor0(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.in_data_reg_88(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.base_address_2(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~0_combout ),
	.base_address_4(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[4]~1_combout ),
	.base_address_3(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~2_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_data_72(\cmd_mux_001|src_data[72]~combout ),
	.src_data_74(\cmd_mux_001|src_data[74]~combout ),
	.src_data_73(\cmd_mux_001|src_data[73]~combout ),
	.src_payload1(\cmd_mux_001|src_payload~1_combout ),
	.src_payload2(\cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\cmd_mux_001|src_payload~3_combout ),
	.src_payload4(\cmd_mux_001|src_payload~4_combout ),
	.src_payload5(\cmd_mux_001|src_payload~5_combout ),
	.src_payload6(\cmd_mux_001|src_payload~6_combout ),
	.src_payload7(\cmd_mux_001|src_payload~7_combout ),
	.src_payload8(\cmd_mux_001|src_payload~8_combout ),
	.src_payload9(\cmd_mux_001|src_payload~9_combout ),
	.src_payload10(\cmd_mux_001|src_payload~10_combout ),
	.src_payload11(\cmd_mux_001|src_payload~11_combout ),
	.src_payload12(\cmd_mux_001|src_payload~12_combout ),
	.src_payload13(\cmd_mux_001|src_payload~13_combout ),
	.src_payload14(\cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\cmd_mux_001|src_payload~15_combout ),
	.src_payload16(\cmd_mux_001|src_payload~16_combout ),
	.src_payload17(\cmd_mux_001|src_payload~17_combout ),
	.src_payload18(\cmd_mux_001|src_payload~18_combout ),
	.src_payload19(\cmd_mux_001|src_payload~19_combout ),
	.src_payload20(\cmd_mux_001|src_payload~20_combout ),
	.src_payload21(\cmd_mux_001|src_payload~21_combout ),
	.src_payload22(\cmd_mux_001|src_payload~22_combout ),
	.src_payload23(\cmd_mux_001|src_payload~23_combout ),
	.src_payload24(\cmd_mux_001|src_payload~24_combout ),
	.src_payload25(\cmd_mux_001|src_payload~25_combout ),
	.src_payload26(\cmd_mux_001|src_payload~26_combout ),
	.src_payload27(\cmd_mux_001|src_payload~27_combout ),
	.src_payload28(\cmd_mux_001|src_payload~28_combout ),
	.src_payload29(\cmd_mux_001|src_payload~29_combout ),
	.src_payload30(\cmd_mux_001|src_payload~30_combout ),
	.src_payload31(\cmd_mux_001|src_payload~31_combout ),
	.src_data_88(\cmd_mux_001|src_data[88]~combout ),
	.src_data_89(\cmd_mux_001|src_data[89]~combout ),
	.src_data_90(\cmd_mux_001|src_data[90]~combout ),
	.src_data_91(\cmd_mux_001|src_data[91]~combout ),
	.src_data_92(\cmd_mux_001|src_data[92]~combout ),
	.src_data_93(\cmd_mux_001|src_data[93]~combout ),
	.src_data_94(\cmd_mux_001|src_data[94]~combout ),
	.src_data_95(\cmd_mux_001|src_data[95]~combout ),
	.src_data_96(\cmd_mux_001|src_data[96]~combout ),
	.src_data_97(\cmd_mux_001|src_data[97]~combout ),
	.src_data_98(\cmd_mux_001|src_data[98]~combout ),
	.src_data_99(\cmd_mux_001|src_data[99]~combout ),
	.src_data_77(\cmd_mux_001|src_data[77]~combout ),
	.out_data_1(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~1_combout ),
	.src_data_71(\cmd_mux_001|src_data[71]~combout ),
	.out_data_0(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~2_combout ),
	.src_data_70(\cmd_mux_001|src_data[70]~combout ));

Computer_System_altera_merlin_burst_adapter dma_1_control_port_slave_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.outclk_wire_0(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.stateST_COMP_TRANS(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(WideOr01),
	.read_latency_shift_reg(\dma_1_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.cp_ready(\dma_1_control_port_slave_agent|cp_ready~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.awready(\arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.r_sync_rst(r_sync_rst),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_59(in_data_reg_59),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.write_cp_data_65(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~0_combout ),
	.write_cp_data_66(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ),
	.write_cp_data_67(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.write_cp_data_68(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ),
	.Add2(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.write_cp_data_69(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~4_combout ),
	.Add21(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.WideNor0(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.nxt_out_eop(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.cmd_src_valid_0(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~2_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.cp_ready1(\dma_1_control_port_slave_agent|cp_ready~2_combout ),
	.in_data_reg_60(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.out_uncomp_byte_cnt_reg_3(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_byte_cnt_reg_2(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_6(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.cmd_src_valid_01(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~3_combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.in_data_reg_88(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_0(in_data_reg_01),
	.in_data_reg_1(in_data_reg_110),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.base_address_2(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~0_combout ),
	.src_data_72(\cmd_mux|src_data[72]~combout ),
	.base_address_4(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[4]~1_combout ),
	.src_data_74(\cmd_mux|src_data[74]~combout ),
	.base_address_3(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~2_combout ),
	.src_data_73(\cmd_mux|src_data[73]~combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.src_payload3(\cmd_mux|src_payload~3_combout ),
	.src_payload4(\cmd_mux|src_payload~4_combout ),
	.src_payload5(\cmd_mux|src_payload~5_combout ),
	.src_payload6(\cmd_mux|src_payload~6_combout ),
	.src_payload7(\cmd_mux|src_payload~7_combout ),
	.src_payload8(\cmd_mux|src_payload~8_combout ),
	.src_payload9(\cmd_mux|src_payload~9_combout ),
	.src_payload10(\cmd_mux|src_payload~10_combout ),
	.src_payload11(\cmd_mux|src_payload~11_combout ),
	.src_payload12(\cmd_mux|src_payload~12_combout ),
	.src_payload13(\cmd_mux|src_payload~13_combout ),
	.src_payload14(\cmd_mux|src_payload~14_combout ),
	.src_payload15(\cmd_mux|src_payload~15_combout ),
	.src_payload16(\cmd_mux|src_payload~16_combout ),
	.src_payload17(\cmd_mux|src_payload~17_combout ),
	.src_payload18(\cmd_mux|src_payload~18_combout ),
	.src_payload19(\cmd_mux|src_payload~19_combout ),
	.src_payload20(\cmd_mux|src_payload~20_combout ),
	.src_payload21(\cmd_mux|src_payload~21_combout ),
	.src_payload22(\cmd_mux|src_payload~22_combout ),
	.src_payload23(\cmd_mux|src_payload~23_combout ),
	.src_payload24(\cmd_mux|src_payload~24_combout ),
	.src_payload25(\cmd_mux|src_payload~25_combout ),
	.src_payload26(\cmd_mux|src_payload~26_combout ),
	.src_payload27(\cmd_mux|src_payload~27_combout ),
	.src_payload28(\cmd_mux|src_payload~28_combout ),
	.src_payload29(\cmd_mux|src_payload~29_combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.src_payload30(\cmd_mux|src_payload~30_combout ),
	.src_payload31(\cmd_mux|src_payload~31_combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.out_data_1(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~1_combout ),
	.src_data_71(\cmd_mux|src_data[71]~combout ),
	.out_data_0(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~2_combout ),
	.src_data_70(\cmd_mux|src_data[70]~combout ));

Computer_System_altera_merlin_traffic_limiter arm_a9_hps_h2f_lw_axi_master_rd_limiter(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_lw_ARADDR_5,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clk(outclk_wire_0),
	.nxt_in_ready(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.WideOr0(\cmd_demux_001|WideOr0~0_combout ),
	.WideOr01(\cmd_demux_001|WideOr0~1_combout ),
	.last_dest_id_0(\arm_a9_hps_h2f_lw_axi_master_rd_limiter|last_dest_id[0]~q ),
	.has_pending_responses1(\arm_a9_hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.cmd_sink_ready(cmd_sink_ready),
	.src1_valid(\rsp_demux|src1_valid~0_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.src1_valid1(\rsp_demux_001|src1_valid~0_combout ),
	.mem_113_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][113]~q ),
	.last_packet_beat(\dma_2_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_channel_0(\arm_a9_hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ),
	.WideOr02(\cmd_demux_001|WideOr0~2_combout ));

Computer_System_altera_merlin_traffic_limiter_1 arm_a9_hps_h2f_lw_axi_master_wr_limiter(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.clk(outclk_wire_0),
	.nxt_in_ready(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.sop_enable(\arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_5(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.WideOr01(\cmd_demux|WideOr0~1_combout ),
	.awready(\arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.src0_valid(\rsp_demux|src0_valid~combout ),
	.src0_valid1(\rsp_demux_001|src0_valid~combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.mem_113_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][113]~q ),
	.last_packet_beat(\dma_2_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.cmd_src_valid_1(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~0_combout ),
	.cmd_src_valid_11(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[1]~1_combout ),
	.cmd_src_valid_0(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~2_combout ),
	.cmd_src_valid_01(\arm_a9_hps_h2f_lw_axi_master_wr_limiter|cmd_src_valid[0]~3_combout ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[5]~0_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.WideOr02(\cmd_demux|WideOr0~2_combout ),
	.WideOr03(\cmd_demux|WideOr0~3_combout ));

Computer_System_altera_avalon_sc_fifo_2 dma_2_control_port_slave_agent_rdata_fifo(
	.clk(outclk_wire_0),
	.read_latency_shift_reg_0(\dma_2_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_2_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\dma_2_control_port_slave_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\dma_2_control_port_slave_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\dma_2_control_port_slave_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\dma_2_control_port_slave_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\dma_2_control_port_slave_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\dma_2_control_port_slave_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\dma_2_control_port_slave_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\dma_2_control_port_slave_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_8(\dma_2_control_port_slave_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_9(\dma_2_control_port_slave_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_10(\dma_2_control_port_slave_translator|av_readdata_pre[10]~q ),
	.mem_10_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_11(\dma_2_control_port_slave_translator|av_readdata_pre[11]~q ),
	.mem_11_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_12(\dma_2_control_port_slave_translator|av_readdata_pre[12]~q ),
	.mem_12_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_13(\dma_2_control_port_slave_translator|av_readdata_pre[13]~q ),
	.mem_13_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_14(\dma_2_control_port_slave_translator|av_readdata_pre[14]~q ),
	.mem_14_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_15(\dma_2_control_port_slave_translator|av_readdata_pre[15]~q ),
	.mem_15_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_16(\dma_2_control_port_slave_translator|av_readdata_pre[16]~q ),
	.mem_16_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_17(\dma_2_control_port_slave_translator|av_readdata_pre[17]~q ),
	.mem_17_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_18(\dma_2_control_port_slave_translator|av_readdata_pre[18]~q ),
	.mem_18_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_19(\dma_2_control_port_slave_translator|av_readdata_pre[19]~q ),
	.mem_19_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_20(\dma_2_control_port_slave_translator|av_readdata_pre[20]~q ),
	.mem_20_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_21(\dma_2_control_port_slave_translator|av_readdata_pre[21]~q ),
	.mem_21_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_22(\dma_2_control_port_slave_translator|av_readdata_pre[22]~q ),
	.mem_22_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_23(\dma_2_control_port_slave_translator|av_readdata_pre[23]~q ),
	.mem_23_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_24(\dma_2_control_port_slave_translator|av_readdata_pre[24]~q ),
	.mem_24_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_25(\dma_2_control_port_slave_translator|av_readdata_pre[25]~q ),
	.mem_25_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_26(\dma_2_control_port_slave_translator|av_readdata_pre[26]~q ),
	.mem_26_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_27(\dma_2_control_port_slave_translator|av_readdata_pre[27]~q ),
	.mem_27_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_28(\dma_2_control_port_slave_translator|av_readdata_pre[28]~q ),
	.mem_28_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_29(\dma_2_control_port_slave_translator|av_readdata_pre[29]~q ),
	.mem_29_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_30(\dma_2_control_port_slave_translator|av_readdata_pre[30]~q ),
	.mem_30_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_31(\dma_2_control_port_slave_translator|av_readdata_pre[31]~q ),
	.mem_31_0(\dma_2_control_port_slave_agent_rdata_fifo|mem[0][31]~q ),
	.reset(r_sync_rst),
	.WideOr0(\rsp_demux_001|WideOr0~0_combout ));

Computer_System_altera_avalon_sc_fifo_3 dma_2_control_port_slave_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.out_valid_reg(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(WideOr0),
	.read_latency_shift_reg(\dma_2_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_112_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_0(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.mem_113_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][113]~q ),
	.comb(\dma_2_control_port_slave_agent|comb~0_combout ),
	.mem_69_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\dma_2_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.mem_88_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][99]~q ),
	.reset(r_sync_rst),
	.in_data_reg_59(in_data_reg_591),
	.mem(mem1),
	.nxt_out_eop(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.WideOr01(\rsp_demux_001|WideOr0~0_combout ),
	.read(\dma_2_control_port_slave_agent_rsp_fifo|read~0_combout ),
	.in_data_reg_60(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.out_uncomp_byte_cnt_reg_6(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_byte_cnt_reg_2(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.rp_valid(\dma_2_control_port_slave_agent|rp_valid~combout ),
	.in_data_reg_88(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ));

Computer_System_altera_merlin_slave_agent_1 dma_2_control_port_slave_agent(
	.outclk_wire_0(outclk_wire_0),
	.stateST_COMP_TRANS(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\dma_2_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(WideOr0),
	.read_latency_shift_reg(\dma_2_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.cp_ready(\dma_2_control_port_slave_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\dma_2_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_2_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\dma_2_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_57_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\dma_2_control_port_slave_agent|comb~0_combout ),
	.mem_69_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\dma_2_control_port_slave_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\dma_2_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.r_sync_rst(r_sync_rst),
	.cp_ready1(\dma_2_control_port_slave_agent|cp_ready~2_combout ),
	.read(\dma_2_control_port_slave_agent_rsp_fifo|read~0_combout ),
	.rp_valid1(\dma_2_control_port_slave_agent|rp_valid~combout ));

Computer_System_altera_avalon_sc_fifo dma_1_control_port_slave_agent_rdata_fifo(
	.clk(outclk_wire_0),
	.read_latency_shift_reg_0(\dma_1_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_1_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\dma_1_control_port_slave_translator|av_readdata_pre[0]~q ),
	.mem_0_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\dma_1_control_port_slave_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\dma_1_control_port_slave_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\dma_1_control_port_slave_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\dma_1_control_port_slave_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\dma_1_control_port_slave_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\dma_1_control_port_slave_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\dma_1_control_port_slave_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_8(\dma_1_control_port_slave_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_9(\dma_1_control_port_slave_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_10(\dma_1_control_port_slave_translator|av_readdata_pre[10]~q ),
	.mem_10_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_11(\dma_1_control_port_slave_translator|av_readdata_pre[11]~q ),
	.mem_11_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_12(\dma_1_control_port_slave_translator|av_readdata_pre[12]~q ),
	.mem_12_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_13(\dma_1_control_port_slave_translator|av_readdata_pre[13]~q ),
	.mem_13_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_14(\dma_1_control_port_slave_translator|av_readdata_pre[14]~q ),
	.mem_14_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_15(\dma_1_control_port_slave_translator|av_readdata_pre[15]~q ),
	.mem_15_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_16(\dma_1_control_port_slave_translator|av_readdata_pre[16]~q ),
	.mem_16_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_17(\dma_1_control_port_slave_translator|av_readdata_pre[17]~q ),
	.mem_17_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_18(\dma_1_control_port_slave_translator|av_readdata_pre[18]~q ),
	.mem_18_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_19(\dma_1_control_port_slave_translator|av_readdata_pre[19]~q ),
	.mem_19_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_20(\dma_1_control_port_slave_translator|av_readdata_pre[20]~q ),
	.mem_20_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_21(\dma_1_control_port_slave_translator|av_readdata_pre[21]~q ),
	.mem_21_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_22(\dma_1_control_port_slave_translator|av_readdata_pre[22]~q ),
	.mem_22_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_23(\dma_1_control_port_slave_translator|av_readdata_pre[23]~q ),
	.mem_23_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_24(\dma_1_control_port_slave_translator|av_readdata_pre[24]~q ),
	.mem_24_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_25(\dma_1_control_port_slave_translator|av_readdata_pre[25]~q ),
	.mem_25_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_26(\dma_1_control_port_slave_translator|av_readdata_pre[26]~q ),
	.mem_26_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_27(\dma_1_control_port_slave_translator|av_readdata_pre[27]~q ),
	.mem_27_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_28(\dma_1_control_port_slave_translator|av_readdata_pre[28]~q ),
	.mem_28_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_29(\dma_1_control_port_slave_translator|av_readdata_pre[29]~q ),
	.mem_29_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_30(\dma_1_control_port_slave_translator|av_readdata_pre[30]~q ),
	.mem_30_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_31(\dma_1_control_port_slave_translator|av_readdata_pre[31]~q ),
	.mem_31_0(\dma_1_control_port_slave_agent_rdata_fifo|mem[0][31]~q ),
	.reset(r_sync_rst),
	.WideOr0(\rsp_demux|WideOr0~0_combout ));

Computer_System_altera_avalon_sc_fifo_1 dma_1_control_port_slave_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.out_valid_reg(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(WideOr01),
	.read_latency_shift_reg(\dma_1_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_112_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_0(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\dma_1_control_port_slave_agent|comb~0_combout ),
	.mem_113_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][113]~q ),
	.mem_65_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][65]~q ),
	.mem_69_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][66]~q ),
	.mem_88_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][99]~q ),
	.reset(r_sync_rst),
	.in_data_reg_59(in_data_reg_59),
	.mem(mem),
	.nxt_out_eop(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.last_packet_beat(\dma_1_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.read(\dma_1_control_port_slave_agent_rsp_fifo|read~0_combout ),
	.in_data_reg_60(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.out_uncomp_byte_cnt_reg_3(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_byte_cnt_reg_2(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_6(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.rp_valid(\dma_1_control_port_slave_agent|rp_valid~combout ),
	.in_data_reg_88(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ));

Computer_System_altera_merlin_slave_agent dma_1_control_port_slave_agent(
	.outclk_wire_0(outclk_wire_0),
	.stateST_COMP_TRANS(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\dma_1_control_port_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(WideOr01),
	.read_latency_shift_reg(\dma_1_control_port_slave_translator|read_latency_shift_reg~0_combout ),
	.cp_ready(\dma_1_control_port_slave_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\dma_1_control_port_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\dma_1_control_port_slave_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\dma_1_control_port_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_57_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\dma_1_control_port_slave_agent|comb~0_combout ),
	.mem_65_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\dma_1_control_port_slave_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\dma_1_control_port_slave_agent_rsp_fifo|mem[0][66]~q ),
	.last_packet_beat1(\dma_1_control_port_slave_agent|uncompressor|last_packet_beat~1_combout ),
	.r_sync_rst(r_sync_rst),
	.cp_ready1(\dma_1_control_port_slave_agent|cp_ready~2_combout ),
	.last_packet_beat2(\dma_1_control_port_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\dma_1_control_port_slave_agent_rsp_fifo|read~0_combout ),
	.rp_valid1(\dma_1_control_port_slave_agent|rp_valid~combout ));

Computer_System_altera_merlin_axi_master_ni arm_a9_hps_h2f_lw_axi_master_agent(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_0(h2f_lw_AWLEN_0),
	.h2f_lw_AWLEN_1(h2f_lw_AWLEN_1),
	.h2f_lw_AWLEN_2(h2f_lw_AWLEN_2),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.outclk_wire_0(outclk_wire_0),
	.sop_enable1(\arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_5(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.awready(\arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.nonposted_cmd_accepted(nonposted_cmd_accepted1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.burst_bytecount_2(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~0_combout ),
	.burst_bytecount_3(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~1_combout ),
	.burst_bytecount_4(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.burst_bytecount_5(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~3_combout ),
	.Add2(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.burst_bytecount_6(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~4_combout ),
	.Add21(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.out_data_5(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[5]~0_combout ),
	.base_address_2(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~0_combout ),
	.Selector4(\arm_a9_hps_h2f_lw_axi_master_agent|Selector4~0_combout ),
	.Selector11(\arm_a9_hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.base_address_4(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[4]~1_combout ),
	.Selector2(\arm_a9_hps_h2f_lw_axi_master_agent|Selector2~0_combout ),
	.Selector9(\arm_a9_hps_h2f_lw_axi_master_agent|Selector9~1_combout ),
	.base_address_3(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~2_combout ),
	.Selector3(\arm_a9_hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\arm_a9_hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.out_data_1(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~1_combout ),
	.Selector5(\arm_a9_hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Selector12(\arm_a9_hps_h2f_lw_axi_master_agent|Selector12~1_combout ),
	.out_data_0(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~2_combout ),
	.Selector6(\arm_a9_hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.Selector13(\arm_a9_hps_h2f_lw_axi_master_agent|Selector13~1_combout ));

endmodule

module Computer_System_altera_avalon_sc_fifo (
	clk,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_9,
	mem_9_0,
	av_readdata_pre_10,
	mem_10_0,
	av_readdata_pre_11,
	mem_11_0,
	av_readdata_pre_12,
	mem_12_0,
	av_readdata_pre_13,
	mem_13_0,
	av_readdata_pre_14,
	mem_14_0,
	av_readdata_pre_15,
	mem_15_0,
	av_readdata_pre_16,
	mem_16_0,
	av_readdata_pre_17,
	mem_17_0,
	av_readdata_pre_18,
	mem_18_0,
	av_readdata_pre_19,
	mem_19_0,
	av_readdata_pre_20,
	mem_20_0,
	av_readdata_pre_21,
	mem_21_0,
	av_readdata_pre_22,
	mem_22_0,
	av_readdata_pre_23,
	mem_23_0,
	av_readdata_pre_24,
	mem_24_0,
	av_readdata_pre_25,
	mem_25_0,
	av_readdata_pre_26,
	mem_26_0,
	av_readdata_pre_27,
	mem_27_0,
	av_readdata_pre_28,
	mem_28_0,
	av_readdata_pre_29,
	mem_29_0,
	av_readdata_pre_30,
	mem_30_0,
	av_readdata_pre_31,
	mem_31_0,
	reset,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	av_readdata_pre_8;
output 	mem_8_0;
input 	av_readdata_pre_9;
output 	mem_9_0;
input 	av_readdata_pre_10;
output 	mem_10_0;
input 	av_readdata_pre_11;
output 	mem_11_0;
input 	av_readdata_pre_12;
output 	mem_12_0;
input 	av_readdata_pre_13;
output 	mem_13_0;
input 	av_readdata_pre_14;
output 	mem_14_0;
input 	av_readdata_pre_15;
output 	mem_15_0;
input 	av_readdata_pre_16;
output 	mem_16_0;
input 	av_readdata_pre_17;
output 	mem_17_0;
input 	av_readdata_pre_18;
output 	mem_18_0;
input 	av_readdata_pre_19;
output 	mem_19_0;
input 	av_readdata_pre_20;
output 	mem_20_0;
input 	av_readdata_pre_21;
output 	mem_21_0;
input 	av_readdata_pre_22;
output 	mem_22_0;
input 	av_readdata_pre_23;
output 	mem_23_0;
input 	av_readdata_pre_24;
output 	mem_24_0;
input 	av_readdata_pre_25;
output 	mem_25_0;
input 	av_readdata_pre_26;
output 	mem_26_0;
input 	av_readdata_pre_27;
output 	mem_27_0;
input 	av_readdata_pre_28;
output 	mem_28_0;
input 	av_readdata_pre_29;
output 	mem_29_0;
input 	av_readdata_pre_30;
output 	mem_30_0;
input 	av_readdata_pre_31;
output 	mem_31_0;
input 	reset;
input 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!av_readdata_pre_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!av_readdata_pre_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!av_readdata_pre_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!av_readdata_pre_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!av_readdata_pre_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!av_readdata_pre_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!av_readdata_pre_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!av_readdata_pre_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!av_readdata_pre_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!av_readdata_pre_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!av_readdata_pre_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!av_readdata_pre_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!av_readdata_pre_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!av_readdata_pre_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!av_readdata_pre_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!av_readdata_pre_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!av_readdata_pre_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!av_readdata_pre_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!av_readdata_pre_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!av_readdata_pre_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!av_readdata_pre_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!av_readdata_pre_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_1 (
	clk,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	read_latency_shift_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_112_0,
	mem_used_0,
	mem_59_0,
	mem_57_0,
	comb,
	mem_113_0,
	mem_65_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	reset,
	in_data_reg_59,
	mem,
	nxt_out_eop,
	last_packet_beat,
	WideOr01,
	read,
	in_data_reg_60,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	rp_valid,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	read_latency_shift_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_112_0;
output 	mem_used_0;
output 	mem_59_0;
output 	mem_57_0;
input 	comb;
output 	mem_113_0;
output 	mem_65_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_88_0;
output 	mem_89_0;
output 	mem_90_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
input 	reset;
input 	in_data_reg_59;
output 	mem;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	WideOr01;
output 	read;
input 	in_data_reg_60;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_6;
input 	rp_valid;
input 	in_data_reg_88;
input 	in_data_reg_89;
input 	in_data_reg_90;
input 	in_data_reg_91;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][112]~q ;
wire \mem~1_combout ;
wire \mem~2_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][59]~q ;
wire \mem~3_combout ;
wire \mem[1][60]~q ;
wire \mem~4_combout ;
wire \mem[1][113]~q ;
wire \mem~5_combout ;
wire \mem[1][65]~q ;
wire \mem~6_combout ;
wire \mem[1][69]~q ;
wire \mem~7_combout ;
wire \mem[1][68]~q ;
wire \mem~8_combout ;
wire \mem[1][67]~q ;
wire \mem~9_combout ;
wire \mem[1][66]~q ;
wire \mem~10_combout ;
wire \mem[1][88]~q ;
wire \mem~11_combout ;
wire \mem[1][89]~q ;
wire \mem~12_combout ;
wire \mem[1][90]~q ;
wire \mem~13_combout ;
wire \mem[1][91]~q ;
wire \mem~14_combout ;
wire \mem[1][92]~q ;
wire \mem~15_combout ;
wire \mem[1][93]~q ;
wire \mem~16_combout ;
wire \mem[1][94]~q ;
wire \mem~17_combout ;
wire \mem[1][95]~q ;
wire \mem~18_combout ;
wire \mem[1][96]~q ;
wire \mem~19_combout ;
wire \mem[1][97]~q ;
wire \mem~20_combout ;
wire \mem[1][98]~q ;
wire \mem~21_combout ;
wire \mem[1][99]~q ;
wire \mem~22_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][88] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_88_0),
	.prn(vcc));
defparam \mem[0][88] .is_wysiwyg = "true";
defparam \mem[0][88] .power_up = "low";

dffeas \mem[0][89] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_89_0),
	.prn(vcc));
defparam \mem[0][89] .is_wysiwyg = "true";
defparam \mem[0][89] .power_up = "low";

dffeas \mem[0][90] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_90_0),
	.prn(vcc));
defparam \mem[0][90] .is_wysiwyg = "true";
defparam \mem[0][90] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4444444444444444;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!WideOr0),
	.datab(!read_latency_shift_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_59),
	.datae(!mem),
	.dataf(!in_data_reg_60),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0000000700007777;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!WideOr0),
	.datab(!nxt_out_eop),
	.datac(!in_data_reg_59),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h0357035703570357;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem~2 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(!\mem[1][112]~q ),
	.datad(!\mem~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0347034703470347;
defparam \mem~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!read),
	.dataf(!\write~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h33331333FFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h2727272727272727;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h2727272727272727;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][113]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h2727272727272727;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h048C37BF048C37BF;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h0437043704370437;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h0437043704370437;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h0437043704370437;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h0437043704370437;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][88] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][88]~q ),
	.prn(vcc));
defparam \mem[1][88] .is_wysiwyg = "true";
defparam \mem[1][88] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][88]~q ),
	.datac(!in_data_reg_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][89]~q ),
	.datac(!in_data_reg_89),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][90] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][90]~q ),
	.prn(vcc));
defparam \mem[1][90] .is_wysiwyg = "true";
defparam \mem[1][90] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][90]~q ),
	.datac(!in_data_reg_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][91]~q ),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~22 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_2 (
	clk,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	av_readdata_pre_0,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_9,
	mem_9_0,
	av_readdata_pre_10,
	mem_10_0,
	av_readdata_pre_11,
	mem_11_0,
	av_readdata_pre_12,
	mem_12_0,
	av_readdata_pre_13,
	mem_13_0,
	av_readdata_pre_14,
	mem_14_0,
	av_readdata_pre_15,
	mem_15_0,
	av_readdata_pre_16,
	mem_16_0,
	av_readdata_pre_17,
	mem_17_0,
	av_readdata_pre_18,
	mem_18_0,
	av_readdata_pre_19,
	mem_19_0,
	av_readdata_pre_20,
	mem_20_0,
	av_readdata_pre_21,
	mem_21_0,
	av_readdata_pre_22,
	mem_22_0,
	av_readdata_pre_23,
	mem_23_0,
	av_readdata_pre_24,
	mem_24_0,
	av_readdata_pre_25,
	mem_25_0,
	av_readdata_pre_26,
	mem_26_0,
	av_readdata_pre_27,
	mem_27_0,
	av_readdata_pre_28,
	mem_28_0,
	av_readdata_pre_29,
	mem_29_0,
	av_readdata_pre_30,
	mem_30_0,
	av_readdata_pre_31,
	mem_31_0,
	reset,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	av_readdata_pre_8;
output 	mem_8_0;
input 	av_readdata_pre_9;
output 	mem_9_0;
input 	av_readdata_pre_10;
output 	mem_10_0;
input 	av_readdata_pre_11;
output 	mem_11_0;
input 	av_readdata_pre_12;
output 	mem_12_0;
input 	av_readdata_pre_13;
output 	mem_13_0;
input 	av_readdata_pre_14;
output 	mem_14_0;
input 	av_readdata_pre_15;
output 	mem_15_0;
input 	av_readdata_pre_16;
output 	mem_16_0;
input 	av_readdata_pre_17;
output 	mem_17_0;
input 	av_readdata_pre_18;
output 	mem_18_0;
input 	av_readdata_pre_19;
output 	mem_19_0;
input 	av_readdata_pre_20;
output 	mem_20_0;
input 	av_readdata_pre_21;
output 	mem_21_0;
input 	av_readdata_pre_22;
output 	mem_22_0;
input 	av_readdata_pre_23;
output 	mem_23_0;
input 	av_readdata_pre_24;
output 	mem_24_0;
input 	av_readdata_pre_25;
output 	mem_25_0;
input 	av_readdata_pre_26;
output 	mem_26_0;
input 	av_readdata_pre_27;
output 	mem_27_0;
input 	av_readdata_pre_28;
output 	mem_28_0;
input 	av_readdata_pre_29;
output 	mem_29_0;
input 	av_readdata_pre_30;
output 	mem_30_0;
input 	av_readdata_pre_31;
output 	mem_31_0;
input 	reset;
input 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!av_readdata_pre_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!av_readdata_pre_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!av_readdata_pre_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!av_readdata_pre_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!av_readdata_pre_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!av_readdata_pre_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!av_readdata_pre_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!av_readdata_pre_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!av_readdata_pre_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!av_readdata_pre_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!av_readdata_pre_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!av_readdata_pre_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!av_readdata_pre_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!av_readdata_pre_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!av_readdata_pre_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!av_readdata_pre_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!av_readdata_pre_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!av_readdata_pre_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!av_readdata_pre_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!av_readdata_pre_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!av_readdata_pre_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!av_readdata_pre_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_3 (
	clk,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	read_latency_shift_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_112_0,
	mem_used_0,
	mem_59_0,
	mem_57_0,
	mem_113_0,
	comb,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	reset,
	in_data_reg_59,
	mem,
	nxt_out_eop,
	WideOr01,
	read,
	in_data_reg_60,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	rp_valid,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	read_latency_shift_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_112_0;
output 	mem_used_0;
output 	mem_59_0;
output 	mem_57_0;
output 	mem_113_0;
input 	comb;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
input 	last_packet_beat;
output 	mem_88_0;
output 	mem_89_0;
output 	mem_90_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
input 	reset;
input 	in_data_reg_59;
output 	mem;
input 	nxt_out_eop;
input 	WideOr01;
output 	read;
input 	in_data_reg_60;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_byte_cnt_reg_2;
input 	rp_valid;
input 	in_data_reg_88;
input 	in_data_reg_89;
input 	in_data_reg_90;
input 	in_data_reg_91;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][112]~q ;
wire \mem~1_combout ;
wire \mem~2_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][59]~q ;
wire \mem~3_combout ;
wire \mem[1][60]~q ;
wire \mem~4_combout ;
wire \mem[1][113]~q ;
wire \mem~5_combout ;
wire \mem[1][69]~q ;
wire \mem~6_combout ;
wire \mem[1][68]~q ;
wire \mem~7_combout ;
wire \mem[1][67]~q ;
wire \mem~8_combout ;
wire \mem[1][66]~q ;
wire \mem~9_combout ;
wire \mem[1][65]~q ;
wire \mem~10_combout ;
wire \mem[1][88]~q ;
wire \mem~11_combout ;
wire \mem[1][89]~q ;
wire \mem~12_combout ;
wire \mem[1][90]~q ;
wire \mem~13_combout ;
wire \mem[1][91]~q ;
wire \mem~14_combout ;
wire \mem[1][92]~q ;
wire \mem~15_combout ;
wire \mem[1][93]~q ;
wire \mem~16_combout ;
wire \mem[1][94]~q ;
wire \mem~17_combout ;
wire \mem[1][95]~q ;
wire \mem~18_combout ;
wire \mem[1][96]~q ;
wire \mem~19_combout ;
wire \mem[1][97]~q ;
wire \mem~20_combout ;
wire \mem[1][98]~q ;
wire \mem~21_combout ;
wire \mem[1][99]~q ;
wire \mem~22_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][88] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_88_0),
	.prn(vcc));
defparam \mem[0][88] .is_wysiwyg = "true";
defparam \mem[0][88] .power_up = "low";

dffeas \mem[0][89] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_89_0),
	.prn(vcc));
defparam \mem[0][89] .is_wysiwyg = "true";
defparam \mem[0][89] .power_up = "low";

dffeas \mem[0][90] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_90_0),
	.prn(vcc));
defparam \mem[0][90] .is_wysiwyg = "true";
defparam \mem[0][90] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4444444444444444;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!WideOr0),
	.datab(!read_latency_shift_reg),
	.datac(!nxt_out_eop),
	.datad(!in_data_reg_59),
	.datae(!mem),
	.dataf(!in_data_reg_60),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0000000700007777;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5505335355053353;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!WideOr0),
	.datab(!nxt_out_eop),
	.datac(!in_data_reg_59),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h0357035703570357;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem~2 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(!\mem[1][112]~q ),
	.datad(!\mem~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0347034703470347;
defparam \mem~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!read),
	.dataf(!\write~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h33331333FFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h2727272727272727;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h2727272727272727;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][113]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h2727272727272727;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0437043704370437;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h0437043704370437;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h0437043704370437;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h0437043704370437;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h048C37BF048C37BF;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][88] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][88]~q ),
	.prn(vcc));
defparam \mem[1][88] .is_wysiwyg = "true";
defparam \mem[1][88] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][88]~q ),
	.datac(!in_data_reg_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][89]~q ),
	.datac(!in_data_reg_89),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][90] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][90]~q ),
	.prn(vcc));
defparam \mem[1][90] .is_wysiwyg = "true";
defparam \mem[1][90] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][90]~q ),
	.datac(!in_data_reg_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][91]~q ),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~22 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_axi_master_ni (
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	outclk_wire_0,
	sop_enable1,
	address_burst_5,
	awready,
	nonposted_cmd_accepted,
	altera_reset_synchronizer_int_chain_out,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_5,
	write_cp_data_68,
	Add2,
	burst_bytecount_6,
	write_cp_data_69,
	Add21,
	out_data_5,
	base_address_2,
	Selector4,
	Selector11,
	base_address_4,
	Selector2,
	Selector9,
	base_address_3,
	Selector3,
	Selector10,
	out_data_1,
	Selector5,
	Selector12,
	out_data_0,
	Selector6,
	Selector13)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	outclk_wire_0;
output 	sop_enable1;
output 	address_burst_5;
output 	awready;
input 	nonposted_cmd_accepted;
input 	altera_reset_synchronizer_int_chain_out;
output 	burst_bytecount_2;
output 	write_cp_data_65;
output 	burst_bytecount_3;
output 	write_cp_data_66;
output 	burst_bytecount_4;
output 	write_cp_data_67;
output 	burst_bytecount_5;
output 	write_cp_data_68;
output 	Add2;
output 	burst_bytecount_6;
output 	write_cp_data_69;
output 	Add21;
output 	out_data_5;
output 	base_address_2;
output 	Selector4;
output 	Selector11;
output 	base_address_4;
output 	Selector2;
output 	Selector9;
output 	base_address_3;
output 	Selector3;
output 	Selector10;
output 	out_data_1;
output 	Selector5;
output 	Selector12;
output 	out_data_0;
output 	Selector6;
output 	Selector13;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|Selector17~0_combout ;
wire \align_address_to_size|Decoder0~1_combout ;
wire \align_address_to_size|Decoder0~2_combout ;
wire \align_address_to_size|Decoder0~3_combout ;
wire \align_address_to_size|Decoder0~4_combout ;
wire \align_address_to_size|Decoder0~5_combout ;
wire \sop_enable~0_combout ;
wire \Add7~0_combout ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add0~0_combout ;
wire \Add7~3_combout ;
wire \log2ceil~0_combout ;
wire \Add1~0_combout ;
wire \Add1~1_combout ;
wire \LessThan12~0_combout ;
wire \Add4~18 ;
wire \Add4~14 ;
wire \Add4~1_sumout ;
wire \Decoder1~0_combout ;
wire \Decoder1~3_combout ;
wire \Decoder1~4_combout ;
wire \Add5~18 ;
wire \Add5~14 ;
wire \Add5~1_sumout ;
wire \log2ceil~1_combout ;
wire \log2ceil~2_combout ;
wire \Selector11~0_combout ;
wire \LessThan14~0_combout ;
wire \Add4~2 ;
wire \Add4~10 ;
wire \Add4~5_sumout ;
wire \Decoder1~1_combout ;
wire \Decoder1~2_combout ;
wire \Add5~2 ;
wire \Add5~10 ;
wire \Add5~5_sumout ;
wire \Selector9~0_combout ;
wire \Add4~9_sumout ;
wire \Add3~0_combout ;
wire \Selector10~0_combout ;
wire \Add5~9_sumout ;
wire \Add4~13_sumout ;
wire \Selector5~0_combout ;
wire \Add5~13_sumout ;
wire \Selector12~0_combout ;
wire \Add4~17_sumout ;
wire \Add5~17_sumout ;
wire \Selector13~0_combout ;


Computer_System_altera_merlin_address_alignment align_address_to_size(
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.clk(outclk_wire_0),
	.sop_enable(sop_enable1),
	.address_burst_5(address_burst_5),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_data_5(out_data_5),
	.log2ceil(\log2ceil~0_combout ),
	.Add1(\Add1~0_combout ),
	.base_address_2(base_address_2),
	.Add11(\Add1~1_combout ),
	.LessThan12(\LessThan12~0_combout ),
	.base_address_4(base_address_4),
	.LessThan14(\LessThan14~0_combout ),
	.base_address_3(base_address_3),
	.Selector17(\align_address_to_size|Selector17~0_combout ),
	.Decoder0(\align_address_to_size|Decoder0~1_combout ),
	.Decoder01(\align_address_to_size|Decoder0~2_combout ),
	.Decoder02(\align_address_to_size|Decoder0~3_combout ),
	.Decoder03(\align_address_to_size|Decoder0~4_combout ),
	.out_data_1(out_data_1),
	.Selector5(\Selector5~0_combout ),
	.Decoder04(\align_address_to_size|Decoder0~5_combout ),
	.out_data_0(out_data_0));

dffeas sop_enable(
	.clk(outclk_wire_0),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

cyclonev_lcell_comb \awready~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(awready),
	.sumout(),
	.cout(),
	.shareout());
defparam \awready~0 .extended_lut = "off";
defparam \awready~0 .lut_mask = 64'h1111111111111111;
defparam \awready~0 .shared_arith = "off";

dffeas \burst_bytecount[2] (
	.clk(outclk_wire_0),
	.d(write_cp_data_65),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_2),
	.prn(vcc));
defparam \burst_bytecount[2] .is_wysiwyg = "true";
defparam \burst_bytecount[2] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[65]~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_65),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[65]~0 .extended_lut = "off";
defparam \write_cp_data[65]~0 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[65]~0 .shared_arith = "off";

dffeas \burst_bytecount[3] (
	.clk(outclk_wire_0),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_3),
	.prn(vcc));
defparam \burst_bytecount[3] .is_wysiwyg = "true";
defparam \burst_bytecount[3] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[66]~1 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[66]~1 .extended_lut = "off";
defparam \write_cp_data[66]~1 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[66]~1 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(outclk_wire_0),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[67]~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[67]~2 .extended_lut = "off";
defparam \write_cp_data[67]~2 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[67]~2 .shared_arith = "off";

dffeas \burst_bytecount[5] (
	.clk(outclk_wire_0),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[68]~3 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_5),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[68]~3 .extended_lut = "off";
defparam \write_cp_data[68]~3 .lut_mask = 64'h478B478B478B478B;
defparam \write_cp_data[68]~3 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add2~0 .shared_arith = "off";

dffeas \burst_bytecount[6] (
	.clk(outclk_wire_0),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_6),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[69]~4 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!\Add0~0_combout ),
	.datad(!burst_bytecount_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[69]~4 .extended_lut = "off";
defparam \write_cp_data[69]~4 .lut_mask = 64'h0437043704370437;
defparam \write_cp_data[69]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0001000100010001;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\LessThan12~0_combout ),
	.datad(!\Add4~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Add5~1_sumout ),
	.datad(!\Selector11~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~1 .extended_lut = "off";
defparam \Selector11~1 .lut_mask = 64'h80A280A280A280A2;
defparam \Selector11~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\LessThan14~0_combout ),
	.datad(!\Add4~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector9~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Add5~5_sumout ),
	.datad(!\Selector9~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector9),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~1 .extended_lut = "off";
defparam \Selector9~1 .lut_mask = 64'h80A280A280A280A2;
defparam \Selector9~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\align_address_to_size|Selector17~0_combout ),
	.datad(!\Add4~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Selector10~0_combout ),
	.datad(!\Add5~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector10~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add4~13_sumout ),
	.datad(!\Selector5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'h80A280A280A280A2;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Add5~13_sumout ),
	.datad(!\Selector12~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~1 .extended_lut = "off";
defparam \Selector12~1 .lut_mask = 64'h80A280A280A280A2;
defparam \Selector12~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add1~1_combout ),
	.datad(!\Add4~17_sumout ),
	.datae(!\Selector5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h8800A8208800A820;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector13~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Decoder1~4_combout ),
	.datad(!\Add5~17_sumout ),
	.datae(!\Selector13~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~1 .extended_lut = "off";
defparam \Selector13~1 .lut_mask = 64'h88008A0288008A02;
defparam \Selector13~1 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_66),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h6666666666666666;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_67),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h4B4B4B4B4B4B4B4B;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_67),
	.datad(!write_cp_data_68),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h40BF40BF40BF40BF;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h0101010101010101;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_67),
	.datad(!write_cp_data_68),
	.datae(!write_cp_data_69),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h4000BFFF4000BFFF;
defparam \Add7~3 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~0 (
	.dataa(!h2f_lw_AWLEN_1),
	.datab(!h2f_lw_AWLEN_2),
	.datac(!h2f_lw_AWLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\log2ceil~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~0 .extended_lut = "off";
defparam \log2ceil~0 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4F00B0FF4F00B0FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan12~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan12~0 .extended_lut = "off";
defparam \LessThan12~0 .lut_mask = 64'hA080800080000000;
defparam \LessThan12~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h00000000000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~17_sumout ),
	.cout(\Add5~18 ),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h00000000000000FF;
defparam \Add5~17 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~13_sumout ),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~1_sumout ),
	.cout(\Add5~2 ),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\log2ceil~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~1 .extended_lut = "off";
defparam \log2ceil~1 .lut_mask = 64'h4F004F004F004F00;
defparam \log2ceil~1 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~2 (
	.dataa(!h2f_lw_ARLEN_1),
	.datab(!h2f_lw_ARLEN_2),
	.datac(!h2f_lw_ARLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\log2ceil~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~2 .extended_lut = "off";
defparam \log2ceil~2 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_0),
	.datac(!h2f_lw_ARSIZE_1),
	.datad(!h2f_lw_ARSIZE_2),
	.datae(!\log2ceil~1_combout ),
	.dataf(!\log2ceil~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'hA800A00080000000;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan14~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan14~0 .extended_lut = "off";
defparam \LessThan14~0 .lut_mask = 64'hE8A0A080A0808000;
defparam \LessThan14~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h0808080808080808;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~9_sumout ),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~5_sumout ),
	.cout(),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_0),
	.datac(!h2f_lw_ARSIZE_1),
	.datad(!h2f_lw_ARSIZE_2),
	.datae(!\log2ceil~1_combout ),
	.dataf(!\log2ceil~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'hEA80AA00A800A000;
defparam \Selector9~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!\Add3~0_combout ),
	.datae(!\log2ceil~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'hA0808000A0808000;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h8000000080000000;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!\Add3~0_combout ),
	.datae(!\log2ceil~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h8000000080000000;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector13~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector13~0 .extended_lut = "off";
defparam \Selector13~0 .lut_mask = 64'h8000800080008000;
defparam \Selector13~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_address_alignment (
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	clk,
	sop_enable,
	address_burst_5,
	nonposted_cmd_accepted,
	reset,
	out_data_5,
	log2ceil,
	Add1,
	base_address_2,
	Add11,
	LessThan12,
	base_address_4,
	LessThan14,
	base_address_3,
	Selector17,
	Decoder0,
	Decoder01,
	Decoder02,
	Decoder03,
	out_data_1,
	Selector5,
	Decoder04,
	out_data_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	clk;
input 	sop_enable;
output 	address_burst_5;
input 	nonposted_cmd_accepted;
input 	reset;
output 	out_data_5;
input 	log2ceil;
input 	Add1;
output 	base_address_2;
input 	Add11;
input 	LessThan12;
output 	base_address_4;
input 	LessThan14;
output 	base_address_3;
output 	Selector17;
output 	Decoder0;
output 	Decoder01;
output 	Decoder02;
output 	Decoder03;
output 	out_data_1;
input 	Selector5;
output 	Decoder04;
output 	out_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~0_combout ;
wire \Add0~21_sumout ;
wire \Add1~21_sumout ;
wire \Selector20~0_combout ;
wire \address_burst[0]~q ;
wire \Add1~22 ;
wire \Add1~17_sumout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \Selector19~0_combout ;
wire \address_burst[1]~q ;
wire \Add1~18 ;
wire \Add1~9_sumout ;
wire \Add0~18 ;
wire \Add0~9_sumout ;
wire \Selector18~0_combout ;
wire \address_burst[2]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Selector17~1_combout ;
wire \address_burst[3]~q ;
wire \Add1~14 ;
wire \Add1~5_sumout ;
wire \Add0~14 ;
wire \Add0~5_sumout ;
wire \Selector16~0_combout ;
wire \address_burst[4]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \address_burst[5]~0_combout ;
wire \address_burst[5]~1_combout ;
wire \address_burst[5]~2_combout ;


dffeas \address_burst[5] (
	.clk(clk),
	.d(\address_burst[5]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(address_burst_5),
	.prn(vcc));
defparam \address_burst[5] .is_wysiwyg = "true";
defparam \address_burst[5] .power_up = "low";

cyclonev_lcell_comb \out_data[5]~0 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~0 .extended_lut = "off";
defparam \out_data[5]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \base_address[2]~0 (
	.dataa(!h2f_lw_AWADDR_2),
	.datab(!sop_enable),
	.datac(!\address_burst[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[2]~0 .extended_lut = "off";
defparam \base_address[2]~0 .lut_mask = 64'h4747474747474747;
defparam \base_address[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \base_address[4]~1 (
	.dataa(!h2f_lw_AWADDR_4),
	.datab(!sop_enable),
	.datac(!\address_burst[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[4]~1 .extended_lut = "off";
defparam \base_address[4]~1 .lut_mask = 64'h4747474747474747;
defparam \base_address[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \base_address[3]~2 (
	.dataa(!h2f_lw_AWADDR_3),
	.datab(!sop_enable),
	.datac(!\address_burst[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[3]~2 .extended_lut = "off";
defparam \base_address[3]~2 .lut_mask = 64'h4747474747474747;
defparam \base_address[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!log2ceil),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector17),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'hA0808000A0808000;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder02),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder03),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~1 (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!sop_enable),
	.datac(!\address_burst[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~1 .extended_lut = "off";
defparam \out_data[1]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder04),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~2 (
	.dataa(!h2f_lw_AWADDR_0),
	.datab(!sop_enable),
	.datac(!\address_burst[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~2 .extended_lut = "off";
defparam \out_data[0]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!sop_enable),
	.datab(!\address_burst[0]~q ),
	.datac(!h2f_lw_AWADDR_0),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!Decoder04),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[0]~q ),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!Add11),
	.datab(!out_data_0),
	.datac(!\Add0~21_sumout ),
	.datad(!\Add1~21_sumout ),
	.datae(!h2f_lw_AWBURST_0),
	.dataf(!h2f_lw_AWBURST_1),
	.datag(!Selector5),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "on";
defparam \Selector20~0 .lut_mask = 64'h33330F0F02F70F0F;
defparam \Selector20~0 .shared_arith = "off";

dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[0]~q ),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add1~17_sumout ),
	.datad(!\Add0~17_sumout ),
	.datae(!out_data_1),
	.dataf(!Selector5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h02578ADF0055AAFF;
defparam \Selector19~0 .shared_arith = "off";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[1]~q ),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!base_address_2),
	.datad(!LessThan12),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector18~0 .shared_arith = "off";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[2]~q ),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Selector17),
	.datad(!base_address_3),
	.datae(!\Add1~13_sumout ),
	.dataf(!\Add0~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~1 .extended_lut = "off";
defparam \Selector17~1 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector17~1 .shared_arith = "off";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector17~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[3]~q ),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!base_address_4),
	.datad(!LessThan14),
	.datae(!\Add1~5_sumout ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector16~0 .shared_arith = "off";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[4]~q ),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_5),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_5),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_5),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_5),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \address_burst[5]~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!log2ceil),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_burst[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_burst[5]~0 .extended_lut = "off";
defparam \address_burst[5]~0 .lut_mask = 64'hE8A0A080E8A0A080;
defparam \address_burst[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \address_burst[5]~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!out_data_5),
	.datad(!\Add1~1_sumout ),
	.datae(!\address_burst[5]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_burst[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_burst[5]~1 .extended_lut = "off";
defparam \address_burst[5]~1 .lut_mask = 64'h082A0A0A082A0A0A;
defparam \address_burst[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \address_burst[5]~2 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!address_burst_5),
	.datac(!nonposted_cmd_accepted),
	.datad(!\Add0~1_sumout ),
	.datae(!\address_burst[5]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_burst[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_burst[5]~2 .extended_lut = "off";
defparam \address_burst[5]~2 .lut_mask = 64'h30353F3F30353F3F;
defparam \address_burst[5]~2 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_adapter (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	outclk_wire_0,
	hold_waitrequest,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	read_latency_shift_reg,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	saved_grant_1,
	saved_grant_0,
	awready,
	r_sync_rst,
	in_data_reg_2,
	in_data_reg_59,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	write_cp_data_65,
	write_cp_data_66,
	write_cp_data_67,
	write_cp_data_68,
	Add2,
	write_cp_data_69,
	Add21,
	WideNor0,
	nxt_out_eop,
	cmd_src_valid_0,
	src0_valid,
	cp_ready1,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	cmd_src_valid_01,
	src_payload_0,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_0,
	in_data_reg_1,
	src_payload,
	base_address_2,
	src_data_72,
	base_address_4,
	src_data_74,
	base_address_3,
	src_data_73,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_payload30,
	src_payload31,
	src_data_77,
	out_data_1,
	src_data_71,
	out_data_0,
	src_data_70)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	outclk_wire_0;
input 	hold_waitrequest;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
input 	mem_used_1;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
input 	read_latency_shift_reg;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	saved_grant_1;
input 	saved_grant_0;
input 	awready;
input 	r_sync_rst;
output 	in_data_reg_2;
output 	in_data_reg_59;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	write_cp_data_65;
input 	write_cp_data_66;
input 	write_cp_data_67;
input 	write_cp_data_68;
input 	Add2;
input 	write_cp_data_69;
input 	Add21;
input 	WideNor0;
output 	nxt_out_eop;
input 	cmd_src_valid_0;
input 	src0_valid;
input 	cp_ready1;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_6;
input 	cmd_src_valid_01;
input 	src_payload_0;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_0;
output 	in_data_reg_1;
input 	src_payload;
input 	base_address_2;
input 	src_data_72;
input 	base_address_4;
input 	src_data_74;
input 	base_address_3;
input 	src_data_73;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_data_88;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_payload30;
input 	src_payload31;
input 	src_data_77;
input 	out_data_1;
input 	src_data_71;
input 	out_data_0;
input 	src_data_70;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_adapter_13_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.outclk_wire_0(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.WideOr01(WideOr0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,src_data_91,src_data_90,src_data_89,src_data_88,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,src_data_77,gnd,gnd,src_data_74,src_data_73,
src_data_72,src_data_71,src_data_70,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,src_payload29,src_payload28,src_payload27,src_payload26,
src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,src_payload6,
src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload,src_payload31,src_payload30}),
	.awready(awready),
	.r_sync_rst(r_sync_rst),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_59(in_data_reg_59),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.write_cp_data_65(write_cp_data_65),
	.write_cp_data_66(write_cp_data_66),
	.write_cp_data_67(write_cp_data_67),
	.write_cp_data_68(write_cp_data_68),
	.Add2(Add2),
	.write_cp_data_69(write_cp_data_69),
	.Add21(Add21),
	.WideNor0(WideNor0),
	.nxt_out_eop(nxt_out_eop),
	.cmd_src_valid_0(cmd_src_valid_0),
	.src0_valid(src0_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_60(in_data_reg_60),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.cmd_src_valid_01(cmd_src_valid_01),
	.sink0_endofpacket(src_payload_0),
	.in_data_reg_88(in_data_reg_88),
	.in_data_reg_89(in_data_reg_89),
	.in_data_reg_90(in_data_reg_90),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.base_address_2(base_address_2),
	.base_address_4(base_address_4),
	.base_address_3(base_address_3),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0));

endmodule

module Computer_System_altera_merlin_burst_adapter_13_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	outclk_wire_0,
	hold_waitrequest,
	stateST_COMP_TRANS,
	out_valid_reg1,
	mem_used_1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr01,
	read_latency_shift_reg,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	sink0_data,
	awready,
	r_sync_rst,
	in_data_reg_2,
	in_data_reg_59,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	write_cp_data_65,
	write_cp_data_66,
	write_cp_data_67,
	write_cp_data_68,
	Add2,
	write_cp_data_69,
	Add21,
	WideNor0,
	nxt_out_eop,
	cmd_src_valid_0,
	src0_valid,
	cp_ready1,
	in_data_reg_60,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	cmd_src_valid_01,
	sink0_endofpacket,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_0,
	in_data_reg_1,
	base_address_2,
	base_address_4,
	base_address_3,
	out_data_1,
	out_data_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	outclk_wire_0;
input 	hold_waitrequest;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
input 	mem_used_1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr01;
input 	read_latency_shift_reg;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	[111:0] sink0_data;
input 	awready;
input 	r_sync_rst;
output 	in_data_reg_2;
output 	in_data_reg_59;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	write_cp_data_65;
input 	write_cp_data_66;
input 	write_cp_data_67;
input 	write_cp_data_68;
input 	Add2;
input 	write_cp_data_69;
input 	Add21;
input 	WideNor0;
output 	nxt_out_eop;
input 	cmd_src_valid_0;
input 	src0_valid;
input 	cp_ready1;
output 	in_data_reg_60;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_6;
input 	cmd_src_valid_01;
input 	sink0_endofpacket;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_0;
output 	in_data_reg_1;
input 	base_address_2;
input 	base_address_4;
input 	base_address_3;
input 	out_data_1;
input 	out_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideOr0~combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \nxt_in_ready~0_combout ;
wire \Selector1~0_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[2]~0_combout ;
wire \d0_int_bytes_remaining[2]~1_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \d0_int_bytes_remaining[3]~2_combout ;
wire \d0_int_bytes_remaining[3]~3_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \d0_int_bytes_remaining[4]~5_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~6_combout ;
wire \d0_int_bytes_remaining[5]~7_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~8_combout ;
wire \d0_int_bytes_remaining[6]~9_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \nxt_in_ready~1_combout ;
wire \nxt_out_eop~0_combout ;
wire \d0_int_nxt_addr[2]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~17_sumout ;
wire \d0_int_nxt_addr[0]~7_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~8_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~6_combout ;
wire \d0_int_nxt_addr[1]~9_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \d0_int_nxt_addr[4]~2_combout ;
wire \in_burstwrap_reg[4]~q ;
wire \nxt_addr[4]~combout ;
wire \int_nxt_addr_reg[4]~q ;
wire \ShiftLeft0~5_combout ;
wire \int_byte_cnt_narrow_reg[4]~0_combout ;
wire \int_byte_cnt_narrow_reg[4]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \Add0~2 ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[4]~3_combout ;
wire \d0_int_nxt_addr[3]~4_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \in_eop_reg~q ;


Computer_System_altera_merlin_address_alignment_1 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_77(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(outclk_wire_0),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(outclk_wire_0),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(outclk_wire_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\nxt_in_ready~1_combout ),
	.datae(gnd),
	.dataf(!\nxt_out_eop~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h11BB11BB10BA10BA;
defparam \nxt_in_ready~2 .shared_arith = "off";

dffeas \in_data_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[59] (
	.clk(outclk_wire_0),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_4),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[4] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(outclk_wire_0),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(outclk_wire_0),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(outclk_wire_0),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(outclk_wire_0),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(outclk_wire_0),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(outclk_wire_0),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(outclk_wire_0),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(outclk_wire_0),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(outclk_wire_0),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(outclk_wire_0),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(outclk_wire_0),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(outclk_wire_0),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(outclk_wire_0),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(outclk_wire_0),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(outclk_wire_0),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(outclk_wire_0),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(outclk_wire_0),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(outclk_wire_0),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(outclk_wire_0),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(outclk_wire_0),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(outclk_wire_0),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(outclk_wire_0),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(outclk_wire_0),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\in_eop_reg~q ),
	.datac(!\nxt_out_eop~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~1 .extended_lut = "off";
defparam \nxt_out_eop~1 .lut_mask = 64'h2727272727272727;
defparam \nxt_out_eop~1 .shared_arith = "off";

dffeas \in_data_reg[60] (
	.clk(outclk_wire_0),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[88] (
	.clk(outclk_wire_0),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_88),
	.prn(vcc));
defparam \in_data_reg[88] .is_wysiwyg = "true";
defparam \in_data_reg[88] .power_up = "low";

dffeas \in_data_reg[89] (
	.clk(outclk_wire_0),
	.d(sink0_data[89]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_89),
	.prn(vcc));
defparam \in_data_reg[89] .is_wysiwyg = "true";
defparam \in_data_reg[89] .power_up = "low";

dffeas \in_data_reg[90] (
	.clk(outclk_wire_0),
	.d(sink0_data[90]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_90),
	.prn(vcc));
defparam \in_data_reg[90] .is_wysiwyg = "true";
defparam \in_data_reg[90] .power_up = "low";

dffeas \in_data_reg[91] (
	.clk(outclk_wire_0),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(outclk_wire_0),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(outclk_wire_0),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(outclk_wire_0),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(outclk_wire_0),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(outclk_wire_0),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(outclk_wire_0),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(outclk_wire_0),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(outclk_wire_0),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!hold_waitrequest),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!awready),
	.datae(!cmd_src_valid_0),
	.dataf(!src0_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000511111115;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!mem_used_1),
	.datac(!WideOr01),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hAEEEAEEEAEEEAEEE;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(outclk_wire_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!nxt_out_eop),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00F800F800F800F8;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!hold_waitrequest),
	.datab(!sink0_data[59]),
	.datac(!cmd_src_valid_01),
	.datad(!\Selector2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0100010001000100;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!out_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h3D3738323D373832;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h10FEBA5410FEBA54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h0D050800F7FFF2FA;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .lut_mask = 64'h1010BA10FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h3D2C3D2C3D2C3D2C;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\WideOr0~combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[60]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h5D55DD5F0C00CC00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\state.ST_IDLE~q ),
	.datab(!\in_valid~combout ),
	.datac(!sink0_data[59]),
	.datad(!nxt_out_eop),
	.datae(!stateST_COMP_TRANS),
	.dataf(!sink0_data[60]),
	.datag(!\nxt_in_ready~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "on";
defparam \Selector1~0 .lut_mask = 64'h0000FF302232FF33;
defparam \Selector1~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~0 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~2 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~2 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~3 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hBF40BF40BF40BF40;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!sink0_data[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'h001E001E001E001E;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[59]),
	.datac(!write_cp_data_67),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~5 .lut_mask = 64'hAB01FF55AB01FF55;
defparam \d0_int_bytes_remaining[4]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4000400040004000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~6 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!write_cp_data_68),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~7 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[6]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~8 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!write_cp_data_69),
	.datad(!Add21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~8 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~9 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~1_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~9 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~9 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~9 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\d0_int_bytes_remaining[2]~1_combout ),
	.datac(!\d0_int_bytes_remaining[3]~3_combout ),
	.datad(!\d0_int_bytes_remaining[4]~5_combout ),
	.datae(!\d0_int_bytes_remaining[5]~7_combout ),
	.dataf(!\d0_int_bytes_remaining[6]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hBAAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(outclk_wire_0),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!nxt_in_ready),
	.datab(!\in_valid~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h2222222222222222;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(outclk_wire_0),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\nxt_in_ready~0_combout ),
	.datab(!nxt_out_eop),
	.datac(!\WideOr0~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h0808080808080808;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!hold_waitrequest),
	.datab(!\nxt_in_ready~0_combout ),
	.datac(!out_valid_reg1),
	.datad(!mem_used_1),
	.datae(!WideOr01),
	.dataf(!read_latency_shift_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h2E2E222E222E222E;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr01),
	.datac(!read_latency_shift_reg),
	.datad(!\new_burst_reg~q ),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_eop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h002AD5FF002AD5FF;
defparam \nxt_out_eop~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~0 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[2]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[72]),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(outclk_wire_0),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~7 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~7 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[0]~q ),
	.datac(!\d0_int_nxt_addr[0]~8_combout ),
	.datad(!sink0_data[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0D080D080D080D08;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~17_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~7_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~8 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~8 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[71]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~6 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~6 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~9 (
	.dataa(!\in_burstwrap_reg[1]~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\int_nxt_addr_reg[1]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(!\d0_int_nxt_addr[1]~6_combout ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~9 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~9 .lut_mask = 64'h1F1F1F1F000000FF;
defparam \d0_int_nxt_addr[1]~9 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[1]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[2]~0_combout ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~2 (
	.dataa(!h2f_lw_ARADDR_4),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~2 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[4]~2 .shared_arith = "off";

dffeas \in_burstwrap_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[74]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[4]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[4] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[4] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[4] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[74]),
	.datac(!\in_burstwrap_reg[4]~q ),
	.datad(!\d0_int_nxt_addr[4]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[4] .extended_lut = "off";
defparam \nxt_addr[4] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[4] .shared_arith = "off";

dffeas \int_nxt_addr_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[4]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!\in_size_reg[0]~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[77]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\new_burst_reg~q ),
	.dataf(!sink0_data[79]),
	.datag(!\in_size_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "on";
defparam \ShiftLeft0~5 .lut_mask = 64'hFF5FFFFFFF5F3F3F;
defparam \ShiftLeft0~5 .shared_arith = "off";

cyclonev_lcell_comb \int_byte_cnt_narrow_reg[4]~0 (
	.dataa(!\ShiftLeft0~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_byte_cnt_narrow_reg[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_byte_cnt_narrow_reg[4]~0 .extended_lut = "off";
defparam \int_byte_cnt_narrow_reg[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \int_byte_cnt_narrow_reg[4]~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[4] (
	.clk(outclk_wire_0),
	.d(\int_byte_cnt_narrow_reg[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[4]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[4] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[4]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[4]~2_combout ),
	.datac(!\int_nxt_addr_reg[4]~q ),
	.datad(!\Add0~5_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~3 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~4 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~4 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[3]~4 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[73]),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[3]~4_combout ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(!\Add0~9_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(outclk_wire_0),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module Computer_System_altera_merlin_address_alignment_1 (
	new_burst_reg,
	src_data_77,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_77;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_77),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_adapter_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	outclk_wire_0,
	hold_waitrequest,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	read_latency_shift_reg,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	saved_grant_1,
	saved_grant_0,
	sop_enable,
	awready,
	r_sync_rst,
	in_data_reg_2,
	in_data_reg_59,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	in_data_reg_0,
	in_data_reg_1,
	nxt_out_eop,
	cmd_src_valid_1,
	src1_valid,
	cp_ready1,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	cmd_src_valid_11,
	src_payload_0,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_5,
	write_cp_data_68,
	Add2,
	burst_bytecount_6,
	write_cp_data_69,
	Add21,
	WideNor0,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	base_address_2,
	base_address_4,
	base_address_3,
	src_payload,
	src_data_72,
	src_data_74,
	src_data_73,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_77,
	out_data_1,
	src_data_71,
	out_data_0,
	src_data_70)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	outclk_wire_0;
input 	hold_waitrequest;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
input 	mem_used_1;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
input 	read_latency_shift_reg;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	saved_grant_1;
input 	saved_grant_0;
input 	sop_enable;
input 	awready;
input 	r_sync_rst;
output 	in_data_reg_2;
output 	in_data_reg_59;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	nxt_out_eop;
input 	cmd_src_valid_1;
input 	src1_valid;
input 	cp_ready1;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_byte_cnt_reg_2;
input 	cmd_src_valid_11;
input 	src_payload_0;
input 	burst_bytecount_2;
input 	write_cp_data_65;
input 	burst_bytecount_3;
input 	write_cp_data_66;
input 	burst_bytecount_4;
input 	write_cp_data_67;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	Add2;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	Add21;
output 	WideNor0;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
input 	base_address_2;
input 	base_address_4;
input 	base_address_3;
input 	src_payload;
input 	src_data_72;
input 	src_data_74;
input 	src_data_73;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_data_88;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_77;
input 	out_data_1;
input 	src_data_71;
input 	out_data_0;
input 	src_data_70;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_adapter_13_1_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.outclk_wire_0(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.WideOr01(WideOr0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.cp_ready(cp_ready),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready(nxt_in_ready),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,src_data_91,src_data_90,src_data_89,src_data_88,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,src_data_77,gnd,gnd,src_data_74,src_data_73,
src_data_72,src_data_71,src_data_70,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,src_payload29,src_payload28,src_payload27,src_payload26,
src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,src_payload6,
src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload,src_payload31,src_payload30}),
	.sop_enable(sop_enable),
	.awready(awready),
	.r_sync_rst(r_sync_rst),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_59(in_data_reg_59),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.nxt_out_eop(nxt_out_eop),
	.cmd_src_valid_1(cmd_src_valid_1),
	.src1_valid(src1_valid),
	.cp_ready1(cp_ready1),
	.in_data_reg_60(in_data_reg_60),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cmd_src_valid_11(cmd_src_valid_11),
	.sink0_endofpacket(src_payload_0),
	.burst_bytecount_2(burst_bytecount_2),
	.write_cp_data_65(write_cp_data_65),
	.burst_bytecount_3(burst_bytecount_3),
	.write_cp_data_66(write_cp_data_66),
	.burst_bytecount_4(burst_bytecount_4),
	.write_cp_data_67(write_cp_data_67),
	.burst_bytecount_5(burst_bytecount_5),
	.write_cp_data_68(write_cp_data_68),
	.Add2(Add2),
	.burst_bytecount_6(burst_bytecount_6),
	.write_cp_data_69(write_cp_data_69),
	.Add21(Add21),
	.WideNor0(WideNor0),
	.in_data_reg_88(in_data_reg_88),
	.in_data_reg_89(in_data_reg_89),
	.in_data_reg_90(in_data_reg_90),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.base_address_2(base_address_2),
	.base_address_4(base_address_4),
	.base_address_3(base_address_3),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0));

endmodule

module Computer_System_altera_merlin_burst_adapter_13_1_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	outclk_wire_0,
	hold_waitrequest,
	stateST_COMP_TRANS,
	out_valid_reg1,
	mem_used_1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr01,
	read_latency_shift_reg,
	cp_ready,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready,
	sink0_data,
	sop_enable,
	awready,
	r_sync_rst,
	in_data_reg_2,
	in_data_reg_59,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	in_data_reg_0,
	in_data_reg_1,
	nxt_out_eop,
	cmd_src_valid_1,
	src1_valid,
	cp_ready1,
	in_data_reg_60,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	cmd_src_valid_11,
	sink0_endofpacket,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_5,
	write_cp_data_68,
	Add2,
	burst_bytecount_6,
	write_cp_data_69,
	Add21,
	WideNor0,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	base_address_2,
	base_address_4,
	base_address_3,
	out_data_1,
	out_data_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	outclk_wire_0;
input 	hold_waitrequest;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
input 	mem_used_1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr01;
input 	read_latency_shift_reg;
input 	cp_ready;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready;
input 	[111:0] sink0_data;
input 	sop_enable;
input 	awready;
input 	r_sync_rst;
output 	in_data_reg_2;
output 	in_data_reg_59;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	nxt_out_eop;
input 	cmd_src_valid_1;
input 	src1_valid;
input 	cp_ready1;
output 	in_data_reg_60;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_byte_cnt_reg_2;
input 	cmd_src_valid_11;
input 	sink0_endofpacket;
input 	burst_bytecount_2;
input 	write_cp_data_65;
input 	burst_bytecount_3;
input 	write_cp_data_66;
input 	burst_bytecount_4;
input 	write_cp_data_67;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	Add2;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	Add21;
output 	WideNor0;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
input 	base_address_2;
input 	base_address_4;
input 	base_address_3;
input 	out_data_1;
input 	out_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideOr0~combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \nxt_in_ready~0_combout ;
wire \Selector1~0_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[2]~0_combout ;
wire \d0_int_bytes_remaining[2]~1_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \d0_int_bytes_remaining[3]~2_combout ;
wire \d0_int_bytes_remaining[3]~3_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \d0_int_bytes_remaining[4]~5_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~6_combout ;
wire \d0_int_bytes_remaining[5]~7_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~8_combout ;
wire \d0_int_bytes_remaining[6]~9_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \nxt_in_ready~1_combout ;
wire \nxt_out_eop~0_combout ;
wire \d0_int_nxt_addr[2]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~17_sumout ;
wire \d0_int_nxt_addr[0]~7_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~8_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~6_combout ;
wire \d0_int_nxt_addr[1]~9_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \d0_int_nxt_addr[4]~2_combout ;
wire \in_burstwrap_reg[4]~q ;
wire \nxt_addr[4]~combout ;
wire \int_nxt_addr_reg[4]~q ;
wire \ShiftLeft0~5_combout ;
wire \int_byte_cnt_narrow_reg[4]~0_combout ;
wire \int_byte_cnt_narrow_reg[4]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \Add0~2 ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[4]~3_combout ;
wire \d0_int_nxt_addr[3]~4_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[3]~5_combout ;
wire \in_eop_reg~q ;


Computer_System_altera_merlin_address_alignment_2 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_77(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(outclk_wire_0),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(outclk_wire_0),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(outclk_wire_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!cp_ready),
	.datad(!\nxt_in_ready~1_combout ),
	.datae(gnd),
	.dataf(!\nxt_out_eop~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h11BB11BB10BA10BA;
defparam \nxt_in_ready~2 .shared_arith = "off";

dffeas \in_data_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[59] (
	.clk(outclk_wire_0),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_4),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[4] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(outclk_wire_0),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(outclk_wire_0),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(outclk_wire_0),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(outclk_wire_0),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(outclk_wire_0),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(outclk_wire_0),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(outclk_wire_0),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(outclk_wire_0),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(outclk_wire_0),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(outclk_wire_0),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(outclk_wire_0),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(outclk_wire_0),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(outclk_wire_0),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(outclk_wire_0),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(outclk_wire_0),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(outclk_wire_0),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(outclk_wire_0),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(outclk_wire_0),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(outclk_wire_0),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(outclk_wire_0),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(outclk_wire_0),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(outclk_wire_0),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(outclk_wire_0),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

dffeas \in_data_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\in_eop_reg~q ),
	.datac(!\nxt_out_eop~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~1 .extended_lut = "off";
defparam \nxt_out_eop~1 .lut_mask = 64'h2727272727272727;
defparam \nxt_out_eop~1 .shared_arith = "off";

dffeas \in_data_reg[60] (
	.clk(outclk_wire_0),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sop_enable),
	.datab(!burst_bytecount_2),
	.datac(!burst_bytecount_3),
	.datad(!burst_bytecount_4),
	.datae(!burst_bytecount_5),
	.dataf(!burst_bytecount_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideNor0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h4000000000000000;
defparam \WideNor0~0 .shared_arith = "off";

dffeas \in_data_reg[88] (
	.clk(outclk_wire_0),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_88),
	.prn(vcc));
defparam \in_data_reg[88] .is_wysiwyg = "true";
defparam \in_data_reg[88] .power_up = "low";

dffeas \in_data_reg[89] (
	.clk(outclk_wire_0),
	.d(sink0_data[89]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_89),
	.prn(vcc));
defparam \in_data_reg[89] .is_wysiwyg = "true";
defparam \in_data_reg[89] .power_up = "low";

dffeas \in_data_reg[90] (
	.clk(outclk_wire_0),
	.d(sink0_data[90]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_90),
	.prn(vcc));
defparam \in_data_reg[90] .is_wysiwyg = "true";
defparam \in_data_reg[90] .power_up = "low";

dffeas \in_data_reg[91] (
	.clk(outclk_wire_0),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(outclk_wire_0),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(outclk_wire_0),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(outclk_wire_0),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(outclk_wire_0),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(outclk_wire_0),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(outclk_wire_0),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(outclk_wire_0),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(outclk_wire_0),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!hold_waitrequest),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!awready),
	.datae(!cmd_src_valid_1),
	.dataf(!src1_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000511111115;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!mem_used_1),
	.datac(!WideOr01),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hAEEEAEEEAEEEAEEE;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(outclk_wire_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!nxt_out_eop),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00F800F800F800F8;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!hold_waitrequest),
	.datab(!sink0_data[59]),
	.datac(!cmd_src_valid_11),
	.datad(!\Selector2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0100010001000100;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_6),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .lut_mask = 64'h337793D733229382;
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_5),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!\Add4~0_combout ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h379D3298379D3298;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_4),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h33D7337733823322;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!out_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .lut_mask = 64'h3D3738323D373832;
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h3D2C3D2C3D2C3D2C;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\Selector2~1_combout ),
	.datab(!\WideOr0~combout ),
	.datac(!\in_valid~combout ),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[60]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h5D55DD5F0C00CC00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\state.ST_IDLE~q ),
	.datab(!\in_valid~combout ),
	.datac(!sink0_data[59]),
	.datad(!nxt_out_eop),
	.datae(!stateST_COMP_TRANS),
	.dataf(!sink0_data[60]),
	.datag(!\nxt_in_ready~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "on";
defparam \Selector1~0 .lut_mask = 64'h0000FF302232FF33;
defparam \Selector1~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~0 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~1 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~2 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~2 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~3 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hBF40BF40BF40BF40;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!sink0_data[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'h001E001E001E001E;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[59]),
	.datac(!\Add1~0_combout ),
	.datad(!write_cp_data_67),
	.datae(!\d0_int_bytes_remaining[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~5 .lut_mask = 64'hA0B1F5F5A0B1F5F5;
defparam \d0_int_bytes_remaining[4]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4000400040004000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~6 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!write_cp_data_68),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~6 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~7 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[6]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~8 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!write_cp_data_69),
	.datad(!Add21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~8 .lut_mask = 64'h0357035703570357;
defparam \d0_int_bytes_remaining[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~9 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~1_combout ),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(!\d0_int_bytes_remaining[6]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~9 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~9 .lut_mask = 64'h08A25DF708A25DF7;
defparam \d0_int_bytes_remaining[6]~9 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\d0_int_bytes_remaining[2]~1_combout ),
	.datac(!\d0_int_bytes_remaining[3]~3_combout ),
	.datad(!\d0_int_bytes_remaining[4]~5_combout ),
	.datae(!\d0_int_bytes_remaining[5]~7_combout ),
	.dataf(!\d0_int_bytes_remaining[6]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hBAAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(outclk_wire_0),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~1 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~1 .extended_lut = "off";
defparam \WideNor0~1 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!nxt_in_ready),
	.datab(!\in_valid~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h2222222222222222;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(outclk_wire_0),
	.d(\WideNor0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\nxt_in_ready~0_combout ),
	.datab(!nxt_out_eop),
	.datac(!\WideOr0~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h0808080808080808;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!hold_waitrequest),
	.datab(!\nxt_in_ready~0_combout ),
	.datac(!out_valid_reg1),
	.datad(!mem_used_1),
	.datae(!WideOr01),
	.dataf(!read_latency_shift_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h2E2E222E222E222E;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr01),
	.datac(!read_latency_shift_reg),
	.datad(!\new_burst_reg~q ),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_eop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h002AD5FF002AD5FF;
defparam \nxt_out_eop~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~0 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[2]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[72]),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(outclk_wire_0),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~7 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~7 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~7 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[0]~q ),
	.datac(!\d0_int_nxt_addr[0]~8_combout ),
	.datad(!sink0_data[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0D080D080D080D08;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~17_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~7_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~8 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~8 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[71]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~6 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~6 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~9 (
	.dataa(!\in_burstwrap_reg[1]~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\int_nxt_addr_reg[1]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(!\d0_int_nxt_addr[1]~6_combout ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~9 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~9 .lut_mask = 64'h1F1F1F1F000000FF;
defparam \d0_int_nxt_addr[1]~9 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[1]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[2]~0_combout ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~2 (
	.dataa(!h2f_lw_ARADDR_4),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~2 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[4]~2 .shared_arith = "off";

dffeas \in_burstwrap_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[74]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[4]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[4] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[4] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[4] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[74]),
	.datac(!\in_burstwrap_reg[4]~q ),
	.datad(!\d0_int_nxt_addr[4]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[4] .extended_lut = "off";
defparam \nxt_addr[4] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[4] .shared_arith = "off";

dffeas \int_nxt_addr_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[4]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!\in_size_reg[0]~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[77]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\new_burst_reg~q ),
	.dataf(!sink0_data[79]),
	.datag(!\in_size_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "on";
defparam \ShiftLeft0~5 .lut_mask = 64'hFF5FFFFFFF5F3F3F;
defparam \ShiftLeft0~5 .shared_arith = "off";

cyclonev_lcell_comb \int_byte_cnt_narrow_reg[4]~0 (
	.dataa(!\ShiftLeft0~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_byte_cnt_narrow_reg[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_byte_cnt_narrow_reg[4]~0 .extended_lut = "off";
defparam \int_byte_cnt_narrow_reg[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \int_byte_cnt_narrow_reg[4]~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[4] (
	.clk(outclk_wire_0),
	.d(\int_byte_cnt_narrow_reg[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[4]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[4] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[4]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[4]~2_combout ),
	.datac(!\int_nxt_addr_reg[4]~q ),
	.datad(!\Add0~5_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~3 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~4 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~4 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[3]~4 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[73]),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[3]~4_combout ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(!\Add0~9_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(outclk_wire_0),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module Computer_System_altera_merlin_address_alignment_2 (
	new_burst_reg,
	src_data_77,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_77;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_77),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_slave_agent (
	outclk_wire_0,
	stateST_COMP_TRANS,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	read_latency_shift_reg,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	mem_57_0,
	comb,
	mem_65_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	last_packet_beat1,
	r_sync_rst,
	cp_ready1,
	last_packet_beat2,
	read,
	rp_valid1)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	read_latency_shift_reg;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	mem_57_0;
output 	comb;
input 	mem_65_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
output 	last_packet_beat1;
input 	r_sync_rst;
output 	cp_ready1;
output 	last_packet_beat2;
input 	read;
output 	rp_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~1_combout ;


Computer_System_altera_merlin_burst_uncompressor uncompressor(
	.clk(outclk_wire_0),
	.mem_57_0(mem_57_0),
	.comb(comb),
	.mem_65_0(mem_65_0),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(r_sync_rst),
	.last_packet_beat2(last_packet_beat2),
	.read(read));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hE000000000000000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!read_latency_shift_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_uncompressor (
	clk,
	mem_57_0,
	comb,
	mem_65_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	mem_57_0;
input 	comb;
input 	mem_65_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h8000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3322322233223222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module Computer_System_altera_merlin_slave_agent_1 (
	outclk_wire_0,
	stateST_COMP_TRANS,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	read_latency_shift_reg,
	cp_ready,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	mem_57_0,
	comb,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	r_sync_rst,
	cp_ready1,
	read,
	rp_valid1)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	stateST_COMP_TRANS;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	read_latency_shift_reg;
output 	cp_ready;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	mem_57_0;
output 	comb;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat;
input 	r_sync_rst;
output 	cp_ready1;
input 	read;
output 	rp_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~1_combout ;


Computer_System_altera_merlin_burst_uncompressor_1 uncompressor(
	.clk(outclk_wire_0),
	.mem_57_0(mem_57_0),
	.comb(comb),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat(last_packet_beat),
	.reset(r_sync_rst),
	.read(read));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hE000000000000000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!read_latency_shift_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~1_combout ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_uncompressor_1 (
	clk,
	mem_57_0,
	comb,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	reset,
	read)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	mem_57_0;
input 	comb;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat;
input 	reset;
input 	read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \last_packet_beat~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \last_packet_beat~1_combout ;


cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!\burst_uncompress_busy~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!\last_packet_beat~0_combout ),
	.dataf(!\last_packet_beat~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3333333222222222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!last_packet_beat),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~0_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_slave_translator (
	clk,
	hold_waitrequest,
	WideOr0,
	wait_latency_counter_1,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	reset,
	in_data_reg_59,
	mem,
	in_data_reg_60,
	av_readdata)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	hold_waitrequest;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	reset;
input 	in_data_reg_59;
input 	mem;
input 	in_data_reg_60;
input 	[31:0] av_readdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter[1]~1_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!hold_waitrequest),
	.datab(!wait_latency_counter_1),
	.datac(!\wait_latency_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0404040404040404;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!WideOr0),
	.datab(!in_data_reg_59),
	.datac(!mem),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'h020A020A020A020A;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[1]~1 (
	.dataa(!hold_waitrequest),
	.datab(!wait_latency_counter_1),
	.datac(!\wait_latency_counter[0]~q ),
	.datad(!\wait_latency_counter[1]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~1 .extended_lut = "off";
defparam \wait_latency_counter[1]~1 .lut_mask = 64'h0051005100510051;
defparam \wait_latency_counter[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~3 (
	.dataa(!\wait_latency_counter[0]~q ),
	.datab(!\wait_latency_counter[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~3 .extended_lut = "off";
defparam \wait_latency_counter~3 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~3 .shared_arith = "off";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_1),
	.datab(!\wait_latency_counter[0]~q ),
	.datac(!\wait_latency_counter[1]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!WideOr0),
	.datab(!read_latency_shift_reg),
	.datac(!mem),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_slave_translator_1 (
	clk,
	hold_waitrequest,
	WideOr0,
	wait_latency_counter_1,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	reset,
	in_data_reg_59,
	mem,
	in_data_reg_60,
	av_readdata)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	hold_waitrequest;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	reset;
input 	in_data_reg_59;
input 	mem;
input 	in_data_reg_60;
input 	[31:0] av_readdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter[0]~1_combout ;
wire \wait_latency_counter~3_combout ;
wire \wait_latency_counter[0]~q ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!hold_waitrequest),
	.datab(!wait_latency_counter_1),
	.datac(!\wait_latency_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0404040404040404;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!WideOr0),
	.datab(!in_data_reg_59),
	.datac(!mem),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h020A020A020A020A;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~1 (
	.dataa(!hold_waitrequest),
	.datab(!wait_latency_counter_1),
	.datac(!\wait_latency_counter[0]~q ),
	.datad(!\wait_latency_counter[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~1 .extended_lut = "off";
defparam \wait_latency_counter[0]~1 .lut_mask = 64'h0051005100510051;
defparam \wait_latency_counter[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~3 (
	.dataa(!\wait_latency_counter[0]~q ),
	.datab(!\wait_latency_counter[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~3 .extended_lut = "off";
defparam \wait_latency_counter~3 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~3 .shared_arith = "off";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_latency_counter[0]~q ),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_1),
	.datab(!\wait_latency_counter[0]~q ),
	.datac(!\wait_latency_counter[0]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!WideOr0),
	.datab(!read_latency_shift_reg),
	.datac(!mem),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_traffic_limiter (
	h2f_lw_ARVALID_0,
	h2f_lw_RREADY_0,
	cmd_sink_data,
	clk,
	nxt_in_ready,
	nxt_in_ready1,
	WideOr0,
	WideOr01,
	last_dest_id_0,
	has_pending_responses1,
	cmd_sink_ready,
	src1_valid,
	src_payload,
	src1_valid1,
	mem_113_0,
	last_packet_beat,
	reset,
	last_channel_0,
	WideOr02)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_RREADY_0;
input 	[117:0] cmd_sink_data;
input 	clk;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	WideOr0;
input 	WideOr01;
output 	last_dest_id_0;
output 	has_pending_responses1;
output 	cmd_sink_ready;
input 	src1_valid;
input 	src_payload;
input 	src1_valid1;
input 	mem_113_0;
input 	last_packet_beat;
input 	reset;
output 	last_channel_0;
input 	WideOr02;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cmd_sink_ready~0_combout ;
wire \save_dest_id~0_combout ;
wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \last_channel[0]~0_combout ;


dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[87]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_dest_id_0),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

cyclonev_lcell_comb \cmd_sink_ready~1 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!WideOr0),
	.datad(!WideOr01),
	.datae(!\cmd_sink_ready~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_sink_ready~1 .extended_lut = "off";
defparam \cmd_sink_ready~1 .lut_mask = 64'h0ACE00000ACE0000;
defparam \cmd_sink_ready~1 .shared_arith = "off";

dffeas \last_channel[0] (
	.clk(clk),
	.d(\last_channel[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

cyclonev_lcell_comb \cmd_sink_ready~0 (
	.dataa(!cmd_sink_data[87]),
	.datab(!last_dest_id_0),
	.datac(!has_pending_responses1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_sink_ready~0 .extended_lut = "off";
defparam \cmd_sink_ready~0 .lut_mask = 64'h0606060606060606;
defparam \cmd_sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!\cmd_sink_ready~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'h4444444444444444;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb response_sink_accepted(
	.dataa(!h2f_lw_RREADY_0),
	.datab(!src1_valid),
	.datac(!src_payload),
	.datad(!src1_valid1),
	.datae(!mem_113_0),
	.dataf(!last_packet_beat),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam response_sink_accepted.extended_lut = "off";
defparam response_sink_accepted.lut_mask = 64'h0404550404040404;
defparam response_sink_accepted.shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!WideOr0),
	.datad(!WideOr01),
	.datae(!\save_dest_id~0_combout ),
	.dataf(!\response_sink_accepted~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h00000ACEFFFFF531;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[1]~q ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6969696969696969;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!WideOr02),
	.datab(!has_pending_responses1),
	.datac(!\save_dest_id~0_combout ),
	.datad(!\pending_response_count[1]~q ),
	.datae(!\pending_response_count[0]~q ),
	.dataf(!\response_sink_accepted~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h3733333333330133;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \last_channel[0]~0 (
	.dataa(!cmd_sink_data[87]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_channel[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_channel[0]~0 .extended_lut = "off";
defparam \last_channel[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_channel[0]~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_traffic_limiter_1 (
	h2f_lw_BREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_AWADDR_5,
	clk,
	nxt_in_ready,
	nxt_in_ready1,
	sop_enable,
	address_burst_5,
	WideOr0,
	WideOr01,
	awready,
	nonposted_cmd_accepted,
	src0_valid,
	src0_valid1,
	src_payload,
	mem_113_0,
	last_packet_beat,
	nonposted_cmd_accepted1,
	reset,
	cmd_src_valid_1,
	cmd_src_valid_11,
	cmd_src_valid_0,
	cmd_src_valid_01,
	cmd_sink_data,
	WideOr02,
	WideOr03)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_AWADDR_5;
input 	clk;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	sop_enable;
input 	address_burst_5;
input 	WideOr0;
input 	WideOr01;
input 	awready;
output 	nonposted_cmd_accepted;
input 	src0_valid;
input 	src0_valid1;
input 	src_payload;
input 	mem_113_0;
input 	last_packet_beat;
output 	nonposted_cmd_accepted1;
input 	reset;
output 	cmd_src_valid_1;
output 	cmd_src_valid_11;
output 	cmd_src_valid_0;
output 	cmd_src_valid_01;
input 	[117:0] cmd_sink_data;
input 	WideOr02;
input 	WideOr03;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \last_dest_id[0]~q ;
wire \pending_response_count[0]~1_combout ;
wire \cmd_sink_ready~0_combout ;
wire \response_sink_accepted~0_combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~q ;
wire \save_dest_id~0_combout ;
wire \last_channel[0]~0_combout ;
wire \last_channel[0]~q ;


cyclonev_lcell_comb \nonposted_cmd_accepted~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(!WideOr0),
	.datae(!WideOr01),
	.dataf(!\save_dest_id~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted),
	.sumout(),
	.cout(),
	.shareout());
defparam \nonposted_cmd_accepted~0 .extended_lut = "off";
defparam \nonposted_cmd_accepted~0 .lut_mask = 64'h0000000000445054;
defparam \nonposted_cmd_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \nonposted_cmd_accepted~1 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!WideOr0),
	.datad(!WideOr01),
	.datae(!\cmd_sink_ready~0_combout ),
	.dataf(!awready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nonposted_cmd_accepted~1 .extended_lut = "off";
defparam \nonposted_cmd_accepted~1 .lut_mask = 64'h000000000ACE0000;
defparam \nonposted_cmd_accepted~1 .shared_arith = "off";

cyclonev_lcell_comb \cmd_src_valid[1]~0 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(!\last_dest_id[0]~q ),
	.datae(!\has_pending_responses~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_src_valid_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_src_valid[1]~0 .extended_lut = "off";
defparam \cmd_src_valid[1]~0 .lut_mask = 64'h4747004747470047;
defparam \cmd_src_valid[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \cmd_src_valid[1]~1 (
	.dataa(!awready),
	.datab(!cmd_src_valid_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_src_valid_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_src_valid[1]~1 .extended_lut = "off";
defparam \cmd_src_valid[1]~1 .lut_mask = 64'h1111111111111111;
defparam \cmd_src_valid[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \cmd_src_valid[0]~2 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(!\has_pending_responses~q ),
	.datae(!\last_channel[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_src_valid_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_src_valid[0]~2 .extended_lut = "off";
defparam \cmd_src_valid[0]~2 .lut_mask = 64'hB800B8B8B800B8B8;
defparam \cmd_src_valid[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \cmd_src_valid[0]~3 (
	.dataa(!awready),
	.datab(!cmd_src_valid_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_src_valid_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_src_valid[0]~3 .extended_lut = "off";
defparam \cmd_src_valid[0]~3 .lut_mask = 64'h1111111111111111;
defparam \cmd_src_valid[0]~3 .shared_arith = "off";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[87]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_dest_id[0]~q ),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \cmd_sink_ready~0 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(!\last_dest_id[0]~q ),
	.datae(!\has_pending_responses~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_sink_ready~0 .extended_lut = "off";
defparam \cmd_sink_ready~0 .lut_mask = 64'h000047B8000047B8;
defparam \cmd_sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!src_payload),
	.datae(!mem_113_0),
	.dataf(!last_packet_beat),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h0011051500110011;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!WideOr02),
	.datac(!WideOr03),
	.datad(!\cmd_sink_ready~0_combout ),
	.datae(!awready),
	.dataf(!\response_sink_accepted~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h00001500FFFFEAFF;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[1]~q ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6969696969696969;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!\has_pending_responses~q ),
	.datab(!nonposted_cmd_accepted),
	.datac(!\pending_response_count[1]~q ),
	.datad(!\pending_response_count[0]~q ),
	.datae(!\response_sink_accepted~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h7555551575555515;
defparam \has_pending_responses~0 .shared_arith = "off";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\has_pending_responses~q ),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(!\last_dest_id[0]~q ),
	.datae(!\has_pending_responses~q ),
	.dataf(!awready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'h00000000FFFFB847;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \last_channel[0]~0 (
	.dataa(!cmd_sink_data[87]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_channel[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_channel[0]~0 .extended_lut = "off";
defparam \last_channel[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_channel[0]~0 .shared_arith = "off";

dffeas \last_channel[0] (
	.clk(clk),
	.d(\last_channel[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(\last_channel[0]~q ),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_demux (
	h2f_lw_AWADDR_5,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_0,
	sop_enable,
	address_burst_5,
	WideOr0,
	saved_grant_01,
	WideOr01,
	WideOr02,
	WideOr03)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_5;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	saved_grant_0;
input 	sop_enable;
input 	address_burst_5;
output 	WideOr0;
input 	saved_grant_01;
output 	WideOr01;
output 	WideOr02;
output 	WideOr03;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!saved_grant_0),
	.datac(!sop_enable),
	.datad(!address_burst_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1013101310131013;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(!saved_grant_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'h00B800B800B800B8;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!nxt_in_ready),
	.datac(!saved_grant_0),
	.datad(!sop_enable),
	.datae(!address_burst_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'h0400040C0400040C;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!nxt_in_ready1),
	.datac(!sop_enable),
	.datad(!address_burst_5),
	.datae(!saved_grant_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr03),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'h00008C8000008C80;
defparam \WideOr0~3 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_demux_1 (
	h2f_lw_ARVALID_0,
	h2f_lw_ARADDR_5,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	WideOr0,
	saved_grant_11,
	WideOr01,
	last_dest_id_0,
	has_pending_responses,
	src1_valid,
	last_channel_0,
	src0_valid,
	WideOr02)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARADDR_5;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	saved_grant_1;
output 	WideOr0;
input 	saved_grant_11;
output 	WideOr01;
input 	last_dest_id_0;
input 	has_pending_responses;
output 	src1_valid;
input 	last_channel_0;
output 	src0_valid;
output 	WideOr02;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_ARADDR_5),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1111111111111111;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!h2f_lw_ARADDR_5),
	.datab(!saved_grant_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'h2222222222222222;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_ARADDR_5),
	.datac(!last_dest_id_0),
	.datad(!has_pending_responses),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h1101110111011101;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_ARADDR_5),
	.datac(!has_pending_responses),
	.datad(!last_channel_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h4044404440444044;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!h2f_lw_ARADDR_5),
	.datab(!saved_grant_1),
	.datac(!nxt_in_ready),
	.datad(!saved_grant_11),
	.datae(!nxt_in_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'h10BA101010BA1010;
defparam \WideOr0~2 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_mux (
	h2f_lw_WLAST_0,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	nxt_in_ready,
	saved_grant_1,
	saved_grant_0,
	awready,
	r_sync_rst,
	cmd_src_valid_0,
	src0_valid,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	cmd_src_valid_01,
	src_payload_0,
	src_payload,
	Selector4,
	Selector11,
	src_data_72,
	Selector2,
	Selector9,
	src_data_74,
	Selector3,
	Selector10,
	src_data_73,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_payload30,
	src_payload31,
	src_data_77,
	Selector5,
	Selector12,
	src_data_71,
	Selector6,
	Selector13,
	src_data_70)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	nxt_in_ready;
output 	saved_grant_1;
output 	saved_grant_0;
input 	awready;
input 	r_sync_rst;
input 	cmd_src_valid_0;
input 	src0_valid;
output 	src_data_78;
output 	src_data_79;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
input 	cmd_src_valid_01;
output 	src_payload_0;
output 	src_payload;
input 	Selector4;
input 	Selector11;
output 	src_data_72;
input 	Selector2;
input 	Selector9;
output 	src_data_74;
input 	Selector3;
input 	Selector10;
output 	src_data_73;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_payload30;
output 	src_payload31;
output 	src_data_77;
input 	Selector5;
input 	Selector12;
output 	src_data_71;
input 	Selector6;
input 	Selector13;
output 	src_data_70;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


Computer_System_altera_merlin_arbitrator_1 arb(
	.clk(outclk_wire_0),
	.nxt_in_ready(nxt_in_ready),
	.reset(r_sync_rst),
	.src0_valid(src0_valid),
	.cmd_src_valid_0(cmd_src_valid_01),
	.src_payload_0(src_payload_0),
	.grant_1(\arb|grant[1]~0_combout ),
	.WideOr1(\WideOr1~combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ));

dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72] .extended_lut = "off";
defparam \src_data[72] .lut_mask = 64'h7530753075307530;
defparam \src_data[72] .shared_arith = "off";

cyclonev_lcell_comb \src_data[74] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector2),
	.datad(!Selector9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74] .extended_lut = "off";
defparam \src_data[74] .lut_mask = 64'h7530753075307530;
defparam \src_data[74] .shared_arith = "off";

cyclonev_lcell_comb \src_data[73] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73] .extended_lut = "off";
defparam \src_data[73] .lut_mask = 64'h7530753075307530;
defparam \src_data[73] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_WDATA_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_WDATA_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_WDATA_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_WDATA_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!h2f_lw_WDATA_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!h2f_lw_WDATA_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!h2f_lw_WDATA_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!h2f_lw_WDATA_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!h2f_lw_WDATA_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!h2f_lw_WDATA_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!h2f_lw_WDATA_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!h2f_lw_WDATA_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!h2f_lw_WDATA_28),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!h2f_lw_WDATA_29),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!h2f_lw_WDATA_30),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!h2f_lw_WDATA_31),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0537053705370537;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0537053705370537;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0537053705370537;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h1111111111111111;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_data[71] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71] .extended_lut = "off";
defparam \src_data[71] .lut_mask = 64'h7530753075307530;
defparam \src_data[71] .shared_arith = "off";

cyclonev_lcell_comb \src_data[70] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70] .extended_lut = "off";
defparam \src_data[70] .lut_mask = 64'h7530753075307530;
defparam \src_data[70] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!awready),
	.datad(!cmd_src_valid_0),
	.datae(!src0_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h0003555700035557;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready),
	.datab(!\WideOr1~combout ),
	.datac(!src_payload_0),
	.datad(!\packet_in_progress~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hCE02CE02CE02CE02;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_mux_1 (
	h2f_lw_WLAST_0,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	nxt_in_ready,
	saved_grant_1,
	saved_grant_0,
	awready,
	r_sync_rst,
	cmd_src_valid_1,
	src1_valid,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	cmd_src_valid_11,
	src_payload_0,
	Selector4,
	Selector11,
	Selector2,
	Selector9,
	Selector3,
	Selector10,
	src_payload,
	src_data_72,
	src_data_74,
	src_data_73,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_77,
	Selector5,
	Selector12,
	src_data_71,
	Selector6,
	Selector13,
	src_data_70)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	nxt_in_ready;
output 	saved_grant_1;
output 	saved_grant_0;
input 	awready;
input 	r_sync_rst;
input 	cmd_src_valid_1;
input 	src1_valid;
output 	src_data_78;
output 	src_data_79;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
input 	cmd_src_valid_11;
output 	src_payload_0;
input 	Selector4;
input 	Selector11;
input 	Selector2;
input 	Selector9;
input 	Selector3;
input 	Selector10;
output 	src_payload;
output 	src_data_72;
output 	src_data_74;
output 	src_data_73;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_77;
input 	Selector5;
input 	Selector12;
output 	src_data_71;
input 	Selector6;
input 	Selector13;
output 	src_data_70;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


Computer_System_altera_merlin_arbitrator arb(
	.clk(outclk_wire_0),
	.nxt_in_ready(nxt_in_ready),
	.reset(r_sync_rst),
	.src1_valid(src1_valid),
	.cmd_src_valid_1(cmd_src_valid_11),
	.src_payload_0(src_payload_0),
	.grant_1(\arb|grant[1]~0_combout ),
	.WideOr1(\WideOr1~combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ));

dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72] .extended_lut = "off";
defparam \src_data[72] .lut_mask = 64'h7530753075307530;
defparam \src_data[72] .shared_arith = "off";

cyclonev_lcell_comb \src_data[74] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector2),
	.datad(!Selector9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74] .extended_lut = "off";
defparam \src_data[74] .lut_mask = 64'h7530753075307530;
defparam \src_data[74] .shared_arith = "off";

cyclonev_lcell_comb \src_data[73] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73] .extended_lut = "off";
defparam \src_data[73] .lut_mask = 64'h7530753075307530;
defparam \src_data[73] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_WDATA_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_WDATA_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_WDATA_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_WDATA_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!h2f_lw_WDATA_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!h2f_lw_WDATA_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!h2f_lw_WDATA_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!h2f_lw_WDATA_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!h2f_lw_WDATA_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!h2f_lw_WDATA_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!h2f_lw_WDATA_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!h2f_lw_WDATA_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!h2f_lw_WDATA_28),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!h2f_lw_WDATA_29),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!h2f_lw_WDATA_30),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!h2f_lw_WDATA_31),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h1111111111111111;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0537053705370537;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0537053705370537;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0537053705370537;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_data[71] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71] .extended_lut = "off";
defparam \src_data[71] .lut_mask = 64'h7530753075307530;
defparam \src_data[71] .shared_arith = "off";

cyclonev_lcell_comb \src_data[70] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!Selector13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70] .extended_lut = "off";
defparam \src_data[70] .lut_mask = 64'h7530753075307530;
defparam \src_data[70] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!awready),
	.datad(!cmd_src_valid_1),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h0003555700035557;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready),
	.datab(!\WideOr1~combout ),
	.datac(!src_payload_0),
	.datad(!\packet_in_progress~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hCE02CE02CE02CE02;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_arbitrator (
	clk,
	nxt_in_ready,
	reset,
	src1_valid,
	cmd_src_valid_1,
	src_payload_0,
	grant_1,
	WideOr1,
	packet_in_progress,
	grant_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	nxt_in_ready;
input 	reset;
input 	src1_valid;
input 	cmd_src_valid_1;
input 	src_payload_0;
output 	grant_1;
input 	WideOr1;
input 	packet_in_progress;
output 	grant_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!cmd_src_valid_1),
	.datad(!src1_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!cmd_src_valid_1),
	.datad(!src1_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!nxt_in_ready),
	.datab(!cmd_src_valid_1),
	.datac(!src1_valid),
	.datad(!WideOr1),
	.datae(!src_payload_0),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h3F003F2A0000002A;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module Computer_System_altera_merlin_arbitrator_1 (
	clk,
	nxt_in_ready,
	reset,
	src0_valid,
	cmd_src_valid_0,
	src_payload_0,
	grant_1,
	WideOr1,
	packet_in_progress,
	grant_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	nxt_in_ready;
input 	reset;
input 	src0_valid;
input 	cmd_src_valid_0;
input 	src_payload_0;
output 	grant_1;
input 	WideOr1;
input 	packet_in_progress;
output 	grant_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!cmd_src_valid_0),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00D500D500D500D5;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!\top_priority_reg[1]~q ),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!cmd_src_valid_0),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0D0C0D0C0D0C0D0C;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!nxt_in_ready),
	.datab(!cmd_src_valid_0),
	.datac(!src0_valid),
	.datad(!WideOr1),
	.datae(!src_payload_0),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h3F003F2A0000002A;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_demux (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_59_0),
	.datad(!mem_57_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_demux_1 (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_59_0),
	.datad(!mem_57_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_mux (
	src0_valid,
	src0_valid1,
	WideOr11,
	mem_88_0,
	mem_88_01,
	src_data_88,
	mem_89_0,
	mem_89_01,
	src_data_89,
	mem_90_0,
	mem_90_01,
	src_data_90,
	mem_91_0,
	mem_91_01,
	src_data_91,
	mem_92_0,
	mem_92_01,
	src_data_92,
	mem_93_0,
	mem_93_01,
	src_data_93,
	mem_94_0,
	mem_94_01,
	src_data_94,
	mem_95_0,
	mem_95_01,
	src_data_95,
	mem_96_0,
	mem_96_01,
	src_data_96,
	mem_97_0,
	mem_97_01,
	src_data_97,
	mem_98_0,
	mem_98_01,
	src_data_98,
	mem_99_0,
	mem_99_01,
	src_data_99)/* synthesis synthesis_greybox=0 */;
input 	src0_valid;
input 	src0_valid1;
output 	WideOr11;
input 	mem_88_0;
input 	mem_88_01;
output 	src_data_88;
input 	mem_89_0;
input 	mem_89_01;
output 	src_data_89;
input 	mem_90_0;
input 	mem_90_01;
output 	src_data_90;
input 	mem_91_0;
input 	mem_91_01;
output 	src_data_91;
input 	mem_92_0;
input 	mem_92_01;
output 	src_data_92;
input 	mem_93_0;
input 	mem_93_01;
output 	src_data_93;
input 	mem_94_0;
input 	mem_94_01;
output 	src_data_94;
input 	mem_95_0;
input 	mem_95_01;
output 	src_data_95;
input 	mem_96_0;
input 	mem_96_01;
output 	src_data_96;
input 	mem_97_0;
input 	mem_97_01;
output 	src_data_97;
input 	mem_98_0;
input 	mem_98_01;
output 	src_data_98;
input 	mem_99_0;
input 	mem_99_01;
output 	src_data_99;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb WideOr1(
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7777777777777777;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_88_0),
	.datad(!mem_88_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_89_0),
	.datad(!mem_89_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0537053705370537;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_90_0),
	.datad(!mem_90_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0537053705370537;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_91_0),
	.datad(!mem_91_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0537053705370537;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_92_0),
	.datad(!mem_92_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_93_0),
	.datad(!mem_93_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_94_0),
	.datad(!mem_94_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_95_0),
	.datad(!mem_95_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_96_0),
	.datad(!mem_96_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_97_0),
	.datad(!mem_97_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_98_0),
	.datad(!mem_98_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!mem_99_0),
	.datad(!mem_99_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_mux_1 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_57_0,
	read_latency_shift_reg_01,
	mem_used_01,
	src1_valid,
	comb,
	mem_113_0,
	mem_65_0,
	last_packet_beat,
	last_packet_beat1,
	src_payload,
	src1_valid1,
	mem_113_01,
	last_packet_beat2,
	src_payload_0,
	WideOr11,
	mem_88_0,
	mem_88_01,
	mem_89_0,
	mem_89_01,
	mem_90_0,
	mem_90_01,
	mem_91_0,
	mem_91_01,
	mem_92_0,
	mem_92_01,
	mem_93_0,
	mem_93_01,
	mem_94_0,
	mem_94_01,
	mem_95_0,
	mem_95_01,
	mem_96_0,
	mem_96_01,
	mem_97_0,
	mem_97_01,
	mem_98_0,
	mem_98_01,
	mem_99_0,
	mem_99_01,
	av_readdata_pre_0,
	mem_0_0,
	av_readdata_pre_01,
	mem_0_01,
	src_data_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_11,
	mem_1_01,
	src_data_1,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_21,
	mem_2_01,
	src_data_2,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_31,
	mem_3_01,
	src_data_3,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_41,
	mem_4_01,
	src_data_4,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_51,
	mem_5_01,
	src_data_5,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_61,
	mem_6_01,
	src_data_6,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_71,
	mem_7_01,
	src_data_7,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_81,
	mem_8_01,
	src_data_8,
	av_readdata_pre_9,
	mem_9_0,
	av_readdata_pre_91,
	mem_9_01,
	src_data_9,
	av_readdata_pre_10,
	mem_10_0,
	av_readdata_pre_101,
	mem_10_01,
	src_data_10,
	av_readdata_pre_111,
	mem_11_0,
	av_readdata_pre_112,
	mem_11_01,
	src_data_11,
	av_readdata_pre_12,
	mem_12_0,
	av_readdata_pre_121,
	mem_12_01,
	src_data_12,
	av_readdata_pre_13,
	mem_13_0,
	av_readdata_pre_131,
	mem_13_01,
	src_data_13,
	av_readdata_pre_14,
	mem_14_0,
	av_readdata_pre_141,
	mem_14_01,
	src_data_14,
	av_readdata_pre_15,
	mem_15_0,
	av_readdata_pre_151,
	mem_15_01,
	src_data_15,
	av_readdata_pre_16,
	mem_16_0,
	av_readdata_pre_161,
	mem_16_01,
	src_data_16,
	av_readdata_pre_17,
	mem_17_0,
	av_readdata_pre_171,
	mem_17_01,
	src_data_17,
	av_readdata_pre_18,
	mem_18_0,
	av_readdata_pre_181,
	mem_18_01,
	src_data_18,
	av_readdata_pre_19,
	mem_19_0,
	av_readdata_pre_191,
	mem_19_01,
	src_data_19,
	av_readdata_pre_20,
	mem_20_0,
	av_readdata_pre_201,
	mem_20_01,
	src_data_20,
	av_readdata_pre_211,
	mem_21_0,
	av_readdata_pre_212,
	mem_21_01,
	src_data_21,
	av_readdata_pre_22,
	mem_22_0,
	av_readdata_pre_221,
	mem_22_01,
	src_data_22,
	av_readdata_pre_23,
	mem_23_0,
	av_readdata_pre_231,
	mem_23_01,
	src_data_23,
	av_readdata_pre_24,
	mem_24_0,
	av_readdata_pre_241,
	mem_24_01,
	src_data_24,
	av_readdata_pre_25,
	mem_25_0,
	av_readdata_pre_251,
	mem_25_01,
	src_data_25,
	av_readdata_pre_26,
	mem_26_0,
	av_readdata_pre_261,
	mem_26_01,
	src_data_26,
	av_readdata_pre_27,
	mem_27_0,
	av_readdata_pre_271,
	mem_27_01,
	src_data_27,
	av_readdata_pre_28,
	mem_28_0,
	av_readdata_pre_281,
	mem_28_01,
	src_data_28,
	av_readdata_pre_29,
	mem_29_0,
	av_readdata_pre_291,
	mem_29_01,
	src_data_29,
	av_readdata_pre_30,
	mem_30_0,
	av_readdata_pre_301,
	mem_30_01,
	src_data_30,
	av_readdata_pre_311,
	mem_31_0,
	av_readdata_pre_312,
	mem_31_01,
	src_data_31,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_57_0;
input 	read_latency_shift_reg_01;
input 	mem_used_01;
input 	src1_valid;
input 	comb;
input 	mem_113_0;
input 	mem_65_0;
input 	last_packet_beat;
input 	last_packet_beat1;
output 	src_payload;
input 	src1_valid1;
input 	mem_113_01;
input 	last_packet_beat2;
output 	src_payload_0;
output 	WideOr11;
input 	mem_88_0;
input 	mem_88_01;
input 	mem_89_0;
input 	mem_89_01;
input 	mem_90_0;
input 	mem_90_01;
input 	mem_91_0;
input 	mem_91_01;
input 	mem_92_0;
input 	mem_92_01;
input 	mem_93_0;
input 	mem_93_01;
input 	mem_94_0;
input 	mem_94_01;
input 	mem_95_0;
input 	mem_95_01;
input 	mem_96_0;
input 	mem_96_01;
input 	mem_97_0;
input 	mem_97_01;
input 	mem_98_0;
input 	mem_98_01;
input 	mem_99_0;
input 	mem_99_01;
input 	av_readdata_pre_0;
input 	mem_0_0;
input 	av_readdata_pre_01;
input 	mem_0_01;
output 	src_data_0;
input 	av_readdata_pre_1;
input 	mem_1_0;
input 	av_readdata_pre_11;
input 	mem_1_01;
output 	src_data_1;
input 	av_readdata_pre_2;
input 	mem_2_0;
input 	av_readdata_pre_21;
input 	mem_2_01;
output 	src_data_2;
input 	av_readdata_pre_3;
input 	mem_3_0;
input 	av_readdata_pre_31;
input 	mem_3_01;
output 	src_data_3;
input 	av_readdata_pre_4;
input 	mem_4_0;
input 	av_readdata_pre_41;
input 	mem_4_01;
output 	src_data_4;
input 	av_readdata_pre_5;
input 	mem_5_0;
input 	av_readdata_pre_51;
input 	mem_5_01;
output 	src_data_5;
input 	av_readdata_pre_6;
input 	mem_6_0;
input 	av_readdata_pre_61;
input 	mem_6_01;
output 	src_data_6;
input 	av_readdata_pre_7;
input 	mem_7_0;
input 	av_readdata_pre_71;
input 	mem_7_01;
output 	src_data_7;
input 	av_readdata_pre_8;
input 	mem_8_0;
input 	av_readdata_pre_81;
input 	mem_8_01;
output 	src_data_8;
input 	av_readdata_pre_9;
input 	mem_9_0;
input 	av_readdata_pre_91;
input 	mem_9_01;
output 	src_data_9;
input 	av_readdata_pre_10;
input 	mem_10_0;
input 	av_readdata_pre_101;
input 	mem_10_01;
output 	src_data_10;
input 	av_readdata_pre_111;
input 	mem_11_0;
input 	av_readdata_pre_112;
input 	mem_11_01;
output 	src_data_11;
input 	av_readdata_pre_12;
input 	mem_12_0;
input 	av_readdata_pre_121;
input 	mem_12_01;
output 	src_data_12;
input 	av_readdata_pre_13;
input 	mem_13_0;
input 	av_readdata_pre_131;
input 	mem_13_01;
output 	src_data_13;
input 	av_readdata_pre_14;
input 	mem_14_0;
input 	av_readdata_pre_141;
input 	mem_14_01;
output 	src_data_14;
input 	av_readdata_pre_15;
input 	mem_15_0;
input 	av_readdata_pre_151;
input 	mem_15_01;
output 	src_data_15;
input 	av_readdata_pre_16;
input 	mem_16_0;
input 	av_readdata_pre_161;
input 	mem_16_01;
output 	src_data_16;
input 	av_readdata_pre_17;
input 	mem_17_0;
input 	av_readdata_pre_171;
input 	mem_17_01;
output 	src_data_17;
input 	av_readdata_pre_18;
input 	mem_18_0;
input 	av_readdata_pre_181;
input 	mem_18_01;
output 	src_data_18;
input 	av_readdata_pre_19;
input 	mem_19_0;
input 	av_readdata_pre_191;
input 	mem_19_01;
output 	src_data_19;
input 	av_readdata_pre_20;
input 	mem_20_0;
input 	av_readdata_pre_201;
input 	mem_20_01;
output 	src_data_20;
input 	av_readdata_pre_211;
input 	mem_21_0;
input 	av_readdata_pre_212;
input 	mem_21_01;
output 	src_data_21;
input 	av_readdata_pre_22;
input 	mem_22_0;
input 	av_readdata_pre_221;
input 	mem_22_01;
output 	src_data_22;
input 	av_readdata_pre_23;
input 	mem_23_0;
input 	av_readdata_pre_231;
input 	mem_23_01;
output 	src_data_23;
input 	av_readdata_pre_24;
input 	mem_24_0;
input 	av_readdata_pre_241;
input 	mem_24_01;
output 	src_data_24;
input 	av_readdata_pre_25;
input 	mem_25_0;
input 	av_readdata_pre_251;
input 	mem_25_01;
output 	src_data_25;
input 	av_readdata_pre_26;
input 	mem_26_0;
input 	av_readdata_pre_261;
input 	mem_26_01;
output 	src_data_26;
input 	av_readdata_pre_27;
input 	mem_27_0;
input 	av_readdata_pre_271;
input 	mem_27_01;
output 	src_data_27;
input 	av_readdata_pre_28;
input 	mem_28_0;
input 	av_readdata_pre_281;
input 	mem_28_01;
output 	src_data_28;
input 	av_readdata_pre_29;
input 	mem_29_0;
input 	av_readdata_pre_291;
input 	mem_29_01;
output 	src_data_29;
input 	av_readdata_pre_30;
input 	mem_30_0;
input 	av_readdata_pre_301;
input 	mem_30_01;
output 	src_data_30;
input 	av_readdata_pre_311;
input 	mem_31_0;
input 	av_readdata_pre_312;
input 	mem_31_01;
output 	src_data_31;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_data[0]~0_combout ;
wire \src_data[0]~1_combout ;
wire \src_data[1]~3_combout ;
wire \src_data[1]~4_combout ;
wire \src_data[2]~6_combout ;
wire \src_data[2]~7_combout ;
wire \src_data[3]~9_combout ;
wire \src_data[3]~10_combout ;
wire \src_data[4]~12_combout ;
wire \src_data[4]~13_combout ;
wire \src_data[5]~15_combout ;
wire \src_data[5]~16_combout ;
wire \src_data[6]~18_combout ;
wire \src_data[6]~19_combout ;
wire \src_data[7]~21_combout ;
wire \src_data[7]~22_combout ;
wire \src_data[8]~24_combout ;
wire \src_data[8]~25_combout ;
wire \src_data[9]~27_combout ;
wire \src_data[9]~28_combout ;
wire \src_data[10]~30_combout ;
wire \src_data[10]~31_combout ;
wire \src_data[11]~33_combout ;
wire \src_data[11]~34_combout ;
wire \src_data[12]~36_combout ;
wire \src_data[12]~37_combout ;
wire \src_data[13]~39_combout ;
wire \src_data[13]~40_combout ;
wire \src_data[14]~42_combout ;
wire \src_data[14]~43_combout ;
wire \src_data[15]~45_combout ;
wire \src_data[15]~46_combout ;
wire \src_data[16]~48_combout ;
wire \src_data[16]~49_combout ;
wire \src_data[17]~51_combout ;
wire \src_data[17]~52_combout ;
wire \src_data[18]~54_combout ;
wire \src_data[18]~55_combout ;
wire \src_data[19]~57_combout ;
wire \src_data[19]~58_combout ;
wire \src_data[20]~60_combout ;
wire \src_data[20]~61_combout ;
wire \src_data[21]~63_combout ;
wire \src_data[21]~64_combout ;
wire \src_data[22]~66_combout ;
wire \src_data[22]~67_combout ;
wire \src_data[23]~69_combout ;
wire \src_data[23]~70_combout ;
wire \src_data[24]~72_combout ;
wire \src_data[24]~73_combout ;
wire \src_data[25]~75_combout ;
wire \src_data[25]~76_combout ;
wire \src_data[26]~78_combout ;
wire \src_data[26]~79_combout ;
wire \src_data[27]~81_combout ;
wire \src_data[27]~82_combout ;
wire \src_data[28]~84_combout ;
wire \src_data[28]~85_combout ;
wire \src_data[29]~87_combout ;
wire \src_data[29]~88_combout ;
wire \src_data[30]~90_combout ;
wire \src_data[30]~91_combout ;
wire \src_data[31]~93_combout ;
wire \src_data[31]~94_combout ;


cyclonev_lcell_comb \src_payload~0 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!mem_113_0),
	.datad(!mem_65_0),
	.datae(!last_packet_beat),
	.dataf(!last_packet_beat1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h0C0C0D0D0C0D0D0D;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!src1_valid),
	.datab(!src_payload),
	.datac(!src1_valid1),
	.datad(!mem_113_01),
	.datae(!last_packet_beat2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h22F2222222F22222;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~2 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[0]~0_combout ),
	.datad(!\src_data[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~2 .extended_lut = "off";
defparam \src_data[0]~2 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~5 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[1]~3_combout ),
	.datad(!\src_data[1]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~5 .extended_lut = "off";
defparam \src_data[1]~5 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~8 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[2]~6_combout ),
	.datad(!\src_data[2]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~8 .extended_lut = "off";
defparam \src_data[2]~8 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[2]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~11 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[3]~9_combout ),
	.datad(!\src_data[3]~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~11 .extended_lut = "off";
defparam \src_data[3]~11 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[3]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~14 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[4]~12_combout ),
	.datad(!\src_data[4]~13_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~14 .extended_lut = "off";
defparam \src_data[4]~14 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[4]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~17 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[5]~15_combout ),
	.datad(!\src_data[5]~16_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~17 .extended_lut = "off";
defparam \src_data[5]~17 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[5]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~20 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[6]~18_combout ),
	.datad(!\src_data[6]~19_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~20 .extended_lut = "off";
defparam \src_data[6]~20 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[6]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~23 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[7]~21_combout ),
	.datad(!\src_data[7]~22_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~23 .extended_lut = "off";
defparam \src_data[7]~23 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[7]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~26 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[8]~24_combout ),
	.datad(!\src_data[8]~25_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~26 .extended_lut = "off";
defparam \src_data[8]~26 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[8]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~29 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[9]~27_combout ),
	.datad(!\src_data[9]~28_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~29 .extended_lut = "off";
defparam \src_data[9]~29 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[9]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~32 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[10]~30_combout ),
	.datad(!\src_data[10]~31_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~32 .extended_lut = "off";
defparam \src_data[10]~32 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[10]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~35 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[11]~33_combout ),
	.datad(!\src_data[11]~34_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~35 .extended_lut = "off";
defparam \src_data[11]~35 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[11]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~38 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[12]~36_combout ),
	.datad(!\src_data[12]~37_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~38 .extended_lut = "off";
defparam \src_data[12]~38 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[12]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~41 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[13]~39_combout ),
	.datad(!\src_data[13]~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~41 .extended_lut = "off";
defparam \src_data[13]~41 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[13]~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~44 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[14]~42_combout ),
	.datad(!\src_data[14]~43_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~44 .extended_lut = "off";
defparam \src_data[14]~44 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[14]~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~47 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[15]~45_combout ),
	.datad(!\src_data[15]~46_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~47 .extended_lut = "off";
defparam \src_data[15]~47 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[15]~47 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~50 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[16]~48_combout ),
	.datad(!\src_data[16]~49_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~50 .extended_lut = "off";
defparam \src_data[16]~50 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[16]~50 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~53 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[17]~51_combout ),
	.datad(!\src_data[17]~52_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~53 .extended_lut = "off";
defparam \src_data[17]~53 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[17]~53 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~56 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[18]~54_combout ),
	.datad(!\src_data[18]~55_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~56 .extended_lut = "off";
defparam \src_data[18]~56 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[18]~56 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~59 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[19]~57_combout ),
	.datad(!\src_data[19]~58_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~59 .extended_lut = "off";
defparam \src_data[19]~59 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[19]~59 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~62 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[20]~60_combout ),
	.datad(!\src_data[20]~61_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~62 .extended_lut = "off";
defparam \src_data[20]~62 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[20]~62 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~65 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[21]~63_combout ),
	.datad(!\src_data[21]~64_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~65 .extended_lut = "off";
defparam \src_data[21]~65 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[21]~65 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~68 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[22]~66_combout ),
	.datad(!\src_data[22]~67_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~68 .extended_lut = "off";
defparam \src_data[22]~68 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[22]~68 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~71 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[23]~69_combout ),
	.datad(!\src_data[23]~70_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~71 .extended_lut = "off";
defparam \src_data[23]~71 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[23]~71 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~74 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[24]~72_combout ),
	.datad(!\src_data[24]~73_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~74 .extended_lut = "off";
defparam \src_data[24]~74 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[24]~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~77 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[25]~75_combout ),
	.datad(!\src_data[25]~76_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~77 .extended_lut = "off";
defparam \src_data[25]~77 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[25]~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~80 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[26]~78_combout ),
	.datad(!\src_data[26]~79_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~80 .extended_lut = "off";
defparam \src_data[26]~80 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[26]~80 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~83 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[27]~81_combout ),
	.datad(!\src_data[27]~82_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~83 .extended_lut = "off";
defparam \src_data[27]~83 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[27]~83 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~86 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[28]~84_combout ),
	.datad(!\src_data[28]~85_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~86 .extended_lut = "off";
defparam \src_data[28]~86 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[28]~86 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~89 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[29]~87_combout ),
	.datad(!\src_data[29]~88_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~89 .extended_lut = "off";
defparam \src_data[29]~89 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[29]~89 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~92 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[30]~90_combout ),
	.datad(!\src_data[30]~91_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~92 .extended_lut = "off";
defparam \src_data[30]~92 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[30]~92 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~95 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!\src_data[31]~93_combout ),
	.datad(!\src_data[31]~94_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~95 .extended_lut = "off";
defparam \src_data[31]~95 .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[31]~95 .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_88_0),
	.datad(!mem_88_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_89_0),
	.datad(!mem_89_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_90_0),
	.datad(!mem_90_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_91_0),
	.datad(!mem_91_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_92_0),
	.datad(!mem_92_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_93_0),
	.datad(!mem_93_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_94_0),
	.datad(!mem_94_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_95_0),
	.datad(!mem_95_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_96_0),
	.datad(!mem_96_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_97_0),
	.datad(!mem_97_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_98_0),
	.datad(!mem_98_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_99_0),
	.datad(!mem_99_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0ACE0ACE0ACE0ACE;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_0),
	.datad(!mem_0_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_01),
	.datad(!mem_0_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_1),
	.datad(!mem_1_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~3 .extended_lut = "off";
defparam \src_data[1]~3 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~4 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_11),
	.datad(!mem_1_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~4 .extended_lut = "off";
defparam \src_data[1]~4 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[1]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~6 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_2),
	.datad(!mem_2_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~6 .extended_lut = "off";
defparam \src_data[2]~6 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~7 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_21),
	.datad(!mem_2_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~7 .extended_lut = "off";
defparam \src_data[2]~7 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[2]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~9 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_3),
	.datad(!mem_3_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~9 .extended_lut = "off";
defparam \src_data[3]~9 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[3]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~10 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_31),
	.datad(!mem_3_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~10 .extended_lut = "off";
defparam \src_data[3]~10 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[3]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~12 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_4),
	.datad(!mem_4_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~12 .extended_lut = "off";
defparam \src_data[4]~12 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[4]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~13 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_41),
	.datad(!mem_4_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~13 .extended_lut = "off";
defparam \src_data[4]~13 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[4]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~15 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_5),
	.datad(!mem_5_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~15 .extended_lut = "off";
defparam \src_data[5]~15 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[5]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~16 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_51),
	.datad(!mem_5_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~16 .extended_lut = "off";
defparam \src_data[5]~16 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[5]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~18 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_6),
	.datad(!mem_6_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~18 .extended_lut = "off";
defparam \src_data[6]~18 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[6]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~19 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_61),
	.datad(!mem_6_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~19 .extended_lut = "off";
defparam \src_data[6]~19 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[6]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~21 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_7),
	.datad(!mem_7_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~21 .extended_lut = "off";
defparam \src_data[7]~21 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[7]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~22 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_71),
	.datad(!mem_7_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~22 .extended_lut = "off";
defparam \src_data[7]~22 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[7]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~24 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_8),
	.datad(!mem_8_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~24 .extended_lut = "off";
defparam \src_data[8]~24 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[8]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~25 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_81),
	.datad(!mem_8_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~25 .extended_lut = "off";
defparam \src_data[8]~25 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[8]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~27 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_9),
	.datad(!mem_9_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~27 .extended_lut = "off";
defparam \src_data[9]~27 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[9]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~28 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_91),
	.datad(!mem_9_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~28 .extended_lut = "off";
defparam \src_data[9]~28 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[9]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~30 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_10),
	.datad(!mem_10_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[10]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~30 .extended_lut = "off";
defparam \src_data[10]~30 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[10]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~31 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_101),
	.datad(!mem_10_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[10]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~31 .extended_lut = "off";
defparam \src_data[10]~31 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[10]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~33 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_111),
	.datad(!mem_11_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[11]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~33 .extended_lut = "off";
defparam \src_data[11]~33 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[11]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~34 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_112),
	.datad(!mem_11_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[11]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~34 .extended_lut = "off";
defparam \src_data[11]~34 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[11]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~36 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_12),
	.datad(!mem_12_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[12]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~36 .extended_lut = "off";
defparam \src_data[12]~36 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[12]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~37 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_121),
	.datad(!mem_12_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[12]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~37 .extended_lut = "off";
defparam \src_data[12]~37 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[12]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~39 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_13),
	.datad(!mem_13_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[13]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~39 .extended_lut = "off";
defparam \src_data[13]~39 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[13]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~40 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_131),
	.datad(!mem_13_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[13]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~40 .extended_lut = "off";
defparam \src_data[13]~40 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[13]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~42 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_14),
	.datad(!mem_14_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[14]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~42 .extended_lut = "off";
defparam \src_data[14]~42 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[14]~42 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~43 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_141),
	.datad(!mem_14_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[14]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~43 .extended_lut = "off";
defparam \src_data[14]~43 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[14]~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~45 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_15),
	.datad(!mem_15_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[15]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~45 .extended_lut = "off";
defparam \src_data[15]~45 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[15]~45 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~46 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_151),
	.datad(!mem_15_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[15]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~46 .extended_lut = "off";
defparam \src_data[15]~46 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[15]~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~48 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_16),
	.datad(!mem_16_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[16]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~48 .extended_lut = "off";
defparam \src_data[16]~48 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[16]~48 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~49 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_161),
	.datad(!mem_16_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[16]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~49 .extended_lut = "off";
defparam \src_data[16]~49 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[16]~49 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~51 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_17),
	.datad(!mem_17_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[17]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~51 .extended_lut = "off";
defparam \src_data[17]~51 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[17]~51 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~52 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_171),
	.datad(!mem_17_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[17]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~52 .extended_lut = "off";
defparam \src_data[17]~52 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[17]~52 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~54 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_18),
	.datad(!mem_18_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[18]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~54 .extended_lut = "off";
defparam \src_data[18]~54 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[18]~54 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~55 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_181),
	.datad(!mem_18_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[18]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~55 .extended_lut = "off";
defparam \src_data[18]~55 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[18]~55 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~57 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_19),
	.datad(!mem_19_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[19]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~57 .extended_lut = "off";
defparam \src_data[19]~57 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[19]~57 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~58 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_191),
	.datad(!mem_19_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[19]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~58 .extended_lut = "off";
defparam \src_data[19]~58 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[19]~58 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~60 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_20),
	.datad(!mem_20_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[20]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~60 .extended_lut = "off";
defparam \src_data[20]~60 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[20]~60 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~61 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_201),
	.datad(!mem_20_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[20]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~61 .extended_lut = "off";
defparam \src_data[20]~61 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[20]~61 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~63 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_211),
	.datad(!mem_21_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[21]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~63 .extended_lut = "off";
defparam \src_data[21]~63 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[21]~63 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~64 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_212),
	.datad(!mem_21_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[21]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~64 .extended_lut = "off";
defparam \src_data[21]~64 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[21]~64 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~66 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_22),
	.datad(!mem_22_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[22]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~66 .extended_lut = "off";
defparam \src_data[22]~66 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[22]~66 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~67 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_221),
	.datad(!mem_22_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[22]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~67 .extended_lut = "off";
defparam \src_data[22]~67 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[22]~67 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~69 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_23),
	.datad(!mem_23_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[23]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~69 .extended_lut = "off";
defparam \src_data[23]~69 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[23]~69 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~70 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_231),
	.datad(!mem_23_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[23]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~70 .extended_lut = "off";
defparam \src_data[23]~70 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[23]~70 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~72 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_24),
	.datad(!mem_24_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[24]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~72 .extended_lut = "off";
defparam \src_data[24]~72 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[24]~72 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~73 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_241),
	.datad(!mem_24_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[24]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~73 .extended_lut = "off";
defparam \src_data[24]~73 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[24]~73 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~75 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_25),
	.datad(!mem_25_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[25]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~75 .extended_lut = "off";
defparam \src_data[25]~75 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[25]~75 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~76 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_251),
	.datad(!mem_25_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[25]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~76 .extended_lut = "off";
defparam \src_data[25]~76 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[25]~76 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~78 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_26),
	.datad(!mem_26_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[26]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~78 .extended_lut = "off";
defparam \src_data[26]~78 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[26]~78 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~79 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_261),
	.datad(!mem_26_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[26]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~79 .extended_lut = "off";
defparam \src_data[26]~79 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[26]~79 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~81 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_27),
	.datad(!mem_27_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~81 .extended_lut = "off";
defparam \src_data[27]~81 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[27]~81 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~82 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_271),
	.datad(!mem_27_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~82 .extended_lut = "off";
defparam \src_data[27]~82 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[27]~82 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~84 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_28),
	.datad(!mem_28_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~84 .extended_lut = "off";
defparam \src_data[28]~84 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[28]~84 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~85 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_281),
	.datad(!mem_28_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~85 .extended_lut = "off";
defparam \src_data[28]~85 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[28]~85 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~87 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_29),
	.datad(!mem_29_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[29]~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~87 .extended_lut = "off";
defparam \src_data[29]~87 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[29]~87 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~88 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_291),
	.datad(!mem_29_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[29]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~88 .extended_lut = "off";
defparam \src_data[29]~88 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[29]~88 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~90 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_30),
	.datad(!mem_30_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~90 .extended_lut = "off";
defparam \src_data[30]~90 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[30]~90 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~91 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_301),
	.datad(!mem_30_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~91 .extended_lut = "off";
defparam \src_data[30]~91 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[30]~91 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~93 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_311),
	.datad(!mem_31_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[31]~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~93 .extended_lut = "off";
defparam \src_data[31]~93 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[31]~93 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~94 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_01),
	.datac(!av_readdata_pre_312),
	.datad(!mem_31_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[31]~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~94 .extended_lut = "off";
defparam \src_data[31]~94 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \src_data[31]~94 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_1 (
	f2h_ARREADY_0,
	f2h_AWREADY_0,
	f2h_BVALID_0,
	f2h_RVALID_0,
	f2h_WREADY_0,
	f2h_RDATA_0,
	f2h_RDATA_1,
	f2h_RDATA_2,
	f2h_RDATA_3,
	f2h_RDATA_4,
	f2h_RDATA_5,
	f2h_RDATA_6,
	f2h_RDATA_7,
	f2h_RDATA_8,
	f2h_RDATA_9,
	f2h_RDATA_10,
	f2h_RDATA_11,
	f2h_RDATA_12,
	f2h_RDATA_13,
	f2h_RDATA_14,
	f2h_RDATA_15,
	f2h_RDATA_16,
	f2h_RDATA_17,
	f2h_RDATA_18,
	f2h_RDATA_19,
	f2h_RDATA_20,
	f2h_RDATA_21,
	f2h_RDATA_22,
	f2h_RDATA_23,
	f2h_RDATA_24,
	f2h_RDATA_25,
	f2h_RDATA_26,
	f2h_RDATA_27,
	f2h_RDATA_28,
	f2h_RDATA_29,
	f2h_RDATA_30,
	f2h_RDATA_31,
	f2h_RDATA_32,
	f2h_RDATA_33,
	f2h_RDATA_34,
	f2h_RDATA_35,
	f2h_RDATA_36,
	f2h_RDATA_37,
	f2h_RDATA_38,
	f2h_RDATA_39,
	f2h_RDATA_40,
	f2h_RDATA_41,
	f2h_RDATA_42,
	f2h_RDATA_43,
	f2h_RDATA_44,
	f2h_RDATA_45,
	f2h_RDATA_46,
	f2h_RDATA_47,
	f2h_RDATA_48,
	f2h_RDATA_49,
	f2h_RDATA_50,
	f2h_RDATA_51,
	f2h_RDATA_52,
	f2h_RDATA_53,
	f2h_RDATA_54,
	f2h_RDATA_55,
	f2h_RDATA_56,
	f2h_RDATA_57,
	f2h_RDATA_58,
	f2h_RDATA_59,
	f2h_RDATA_60,
	f2h_RDATA_61,
	f2h_RDATA_62,
	f2h_RDATA_63,
	outclk_wire_0,
	readaddress_2,
	readaddress_3,
	readaddress_4,
	readaddress_5,
	readaddress_6,
	readaddress_7,
	readaddress_8,
	readaddress_9,
	readaddress_10,
	readaddress_11,
	readaddress_12,
	readaddress_13,
	readaddress_14,
	readaddress_15,
	readaddress_16,
	readaddress_17,
	readaddress_18,
	readaddress_19,
	readaddress_20,
	readaddress_21,
	readaddress_22,
	readaddress_23,
	readaddress_24,
	readaddress_25,
	readaddress_26,
	readaddress_27,
	readaddress_28,
	readaddress_29,
	readaddress_30,
	readaddress_31,
	writeaddress_2,
	writeaddress_3,
	writeaddress_4,
	writeaddress_5,
	writeaddress_6,
	writeaddress_7,
	writeaddress_8,
	writeaddress_9,
	writeaddress_10,
	writeaddress_11,
	writeaddress_12,
	writeaddress_13,
	writeaddress_14,
	writeaddress_15,
	writeaddress_16,
	writeaddress_17,
	writeaddress_18,
	writeaddress_19,
	writeaddress_20,
	writeaddress_21,
	writeaddress_22,
	writeaddress_23,
	writeaddress_24,
	writeaddress_25,
	writeaddress_26,
	writeaddress_27,
	writeaddress_28,
	writeaddress_29,
	writeaddress_30,
	writeaddress_31,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	writeaddress_1,
	writeaddress_0,
	mem_used_7,
	saved_grant_0,
	read_select,
	hold_waitrequest,
	write,
	arvalid,
	address_taken,
	mem_used_71,
	fifo_empty,
	saved_grant_1,
	src_valid,
	awvalid,
	ARM_A9_HPS_f2h_axi_slave_bready,
	data_taken,
	wvalid,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	src_payload50,
	src_payload51,
	src_payload52,
	src_payload53,
	src_payload54,
	src_payload55,
	src_payload56,
	src_payload57,
	src_payload58,
	src_payload59,
	last_write_collision,
	last_write_data_0,
	control_2,
	control_0,
	ShiftLeft1,
	last_write_data_1,
	ShiftLeft11,
	last_write_data_2,
	ShiftLeft12,
	last_write_data_3,
	ShiftLeft13,
	last_write_data_4,
	ShiftLeft14,
	last_write_data_5,
	ShiftLeft15,
	last_write_data_6,
	ShiftLeft16,
	last_write_data_7,
	ShiftLeft17,
	write_writedata,
	last_write_data_8,
	ShiftLeft18,
	write_writedata1,
	last_write_data_9,
	ShiftLeft19,
	write_writedata2,
	last_write_data_10,
	ShiftLeft110,
	write_writedata3,
	last_write_data_11,
	ShiftLeft111,
	write_writedata4,
	last_write_data_12,
	ShiftLeft112,
	write_writedata5,
	last_write_data_13,
	ShiftLeft113,
	write_writedata6,
	last_write_data_14,
	ShiftLeft114,
	write_writedata7,
	last_write_data_15,
	ShiftLeft115,
	last_write_data_16,
	ShiftLeft116,
	last_write_data_17,
	ShiftLeft117,
	last_write_data_18,
	ShiftLeft118,
	last_write_data_19,
	ShiftLeft119,
	last_write_data_20,
	ShiftLeft120,
	last_write_data_21,
	ShiftLeft121,
	last_write_data_22,
	ShiftLeft122,
	last_write_data_23,
	ShiftLeft123,
	last_write_data_24,
	ShiftLeft124,
	last_write_data_25,
	ShiftLeft125,
	last_write_data_26,
	ShiftLeft126,
	last_write_data_27,
	ShiftLeft127,
	last_write_data_28,
	ShiftLeft128,
	last_write_data_29,
	ShiftLeft129,
	last_write_data_30,
	ShiftLeft130,
	last_write_data_31,
	ShiftLeft131,
	ShiftLeft132,
	ShiftLeft133,
	ShiftLeft134,
	ShiftLeft135,
	ShiftLeft136,
	ShiftLeft137,
	ShiftLeft138,
	ShiftLeft139,
	ShiftLeft140,
	ShiftLeft141,
	ShiftLeft142,
	ShiftLeft143,
	ShiftLeft144,
	ShiftLeft145,
	ShiftLeft146,
	ShiftLeft147,
	ShiftLeft148,
	ShiftLeft149,
	ShiftLeft150,
	ShiftLeft151,
	ShiftLeft152,
	ShiftLeft153,
	ShiftLeft154,
	ShiftLeft155,
	ShiftLeft156,
	ShiftLeft157,
	ShiftLeft158,
	ShiftLeft159,
	ShiftLeft160,
	ShiftLeft161,
	ShiftLeft162,
	ShiftLeft163,
	ShiftLeft0,
	ShiftLeft01,
	ShiftLeft02,
	ShiftLeft03,
	ShiftLeft04,
	ShiftLeft05,
	ShiftLeft06,
	ShiftLeft07,
	altera_reset_synchronizer_int_chain_out,
	WideOr1,
	r_sync_rst,
	inc_read,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	av_readdatavalid3,
	fifo_read,
	write_cp_ready,
	av_readdatavalid4,
	src0_valid,
	src_data_8,
	src_data_81,
	src_data_16,
	src_data_24,
	src_data_0,
	src_data_01,
	src_data_9,
	src_data_91,
	src_data_17,
	src_data_25,
	src_data_1,
	src_data_11,
	src_data_10,
	src_data_101,
	src_data_18,
	src_data_26,
	src_data_2,
	src_data_21,
	src_data_111,
	src_data_112,
	src_data_19,
	src_data_27,
	src_data_3,
	src_data_31,
	src_data_12,
	src_data_121,
	src_data_20,
	src_data_28,
	src_data_4,
	src_data_41,
	src_data_13,
	src_data_131,
	src_data_211,
	src_data_29,
	src_data_5,
	src_data_51,
	src_data_14,
	src_data_141,
	src_data_22,
	src_data_30,
	src_data_6,
	src_data_61,
	src_data_15,
	src_data_151,
	src_data_23,
	src_data_311,
	src_data_7,
	src_data_71,
	src_data_82,
	src_data_92,
	src_data_102,
	src_data_113,
	src_data_122,
	src_data_132,
	src_data_142,
	src_data_152)/* synthesis synthesis_greybox=0 */;
input 	f2h_ARREADY_0;
input 	f2h_AWREADY_0;
input 	f2h_BVALID_0;
input 	f2h_RVALID_0;
input 	f2h_WREADY_0;
input 	f2h_RDATA_0;
input 	f2h_RDATA_1;
input 	f2h_RDATA_2;
input 	f2h_RDATA_3;
input 	f2h_RDATA_4;
input 	f2h_RDATA_5;
input 	f2h_RDATA_6;
input 	f2h_RDATA_7;
input 	f2h_RDATA_8;
input 	f2h_RDATA_9;
input 	f2h_RDATA_10;
input 	f2h_RDATA_11;
input 	f2h_RDATA_12;
input 	f2h_RDATA_13;
input 	f2h_RDATA_14;
input 	f2h_RDATA_15;
input 	f2h_RDATA_16;
input 	f2h_RDATA_17;
input 	f2h_RDATA_18;
input 	f2h_RDATA_19;
input 	f2h_RDATA_20;
input 	f2h_RDATA_21;
input 	f2h_RDATA_22;
input 	f2h_RDATA_23;
input 	f2h_RDATA_24;
input 	f2h_RDATA_25;
input 	f2h_RDATA_26;
input 	f2h_RDATA_27;
input 	f2h_RDATA_28;
input 	f2h_RDATA_29;
input 	f2h_RDATA_30;
input 	f2h_RDATA_31;
input 	f2h_RDATA_32;
input 	f2h_RDATA_33;
input 	f2h_RDATA_34;
input 	f2h_RDATA_35;
input 	f2h_RDATA_36;
input 	f2h_RDATA_37;
input 	f2h_RDATA_38;
input 	f2h_RDATA_39;
input 	f2h_RDATA_40;
input 	f2h_RDATA_41;
input 	f2h_RDATA_42;
input 	f2h_RDATA_43;
input 	f2h_RDATA_44;
input 	f2h_RDATA_45;
input 	f2h_RDATA_46;
input 	f2h_RDATA_47;
input 	f2h_RDATA_48;
input 	f2h_RDATA_49;
input 	f2h_RDATA_50;
input 	f2h_RDATA_51;
input 	f2h_RDATA_52;
input 	f2h_RDATA_53;
input 	f2h_RDATA_54;
input 	f2h_RDATA_55;
input 	f2h_RDATA_56;
input 	f2h_RDATA_57;
input 	f2h_RDATA_58;
input 	f2h_RDATA_59;
input 	f2h_RDATA_60;
input 	f2h_RDATA_61;
input 	f2h_RDATA_62;
input 	f2h_RDATA_63;
input 	outclk_wire_0;
input 	readaddress_2;
input 	readaddress_3;
input 	readaddress_4;
input 	readaddress_5;
input 	readaddress_6;
input 	readaddress_7;
input 	readaddress_8;
input 	readaddress_9;
input 	readaddress_10;
input 	readaddress_11;
input 	readaddress_12;
input 	readaddress_13;
input 	readaddress_14;
input 	readaddress_15;
input 	readaddress_16;
input 	readaddress_17;
input 	readaddress_18;
input 	readaddress_19;
input 	readaddress_20;
input 	readaddress_21;
input 	readaddress_22;
input 	readaddress_23;
input 	readaddress_24;
input 	readaddress_25;
input 	readaddress_26;
input 	readaddress_27;
input 	readaddress_28;
input 	readaddress_29;
input 	readaddress_30;
input 	readaddress_31;
input 	writeaddress_2;
input 	writeaddress_3;
input 	writeaddress_4;
input 	writeaddress_5;
input 	writeaddress_6;
input 	writeaddress_7;
input 	writeaddress_8;
input 	writeaddress_9;
input 	writeaddress_10;
input 	writeaddress_11;
input 	writeaddress_12;
input 	writeaddress_13;
input 	writeaddress_14;
input 	writeaddress_15;
input 	writeaddress_16;
input 	writeaddress_17;
input 	writeaddress_18;
input 	writeaddress_19;
input 	writeaddress_20;
input 	writeaddress_21;
input 	writeaddress_22;
input 	writeaddress_23;
input 	writeaddress_24;
input 	writeaddress_25;
input 	writeaddress_26;
input 	writeaddress_27;
input 	writeaddress_28;
input 	writeaddress_29;
input 	writeaddress_30;
input 	writeaddress_31;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	writeaddress_1;
input 	writeaddress_0;
output 	mem_used_7;
output 	saved_grant_0;
input 	read_select;
input 	hold_waitrequest;
output 	write;
output 	arvalid;
output 	address_taken;
output 	mem_used_71;
input 	fifo_empty;
output 	saved_grant_1;
output 	src_valid;
output 	awvalid;
output 	ARM_A9_HPS_f2h_axi_slave_bready;
output 	data_taken;
output 	wvalid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
output 	src_payload35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	src_payload46;
output 	src_payload47;
output 	src_payload48;
output 	src_payload49;
output 	src_payload50;
output 	src_payload51;
output 	src_payload52;
output 	src_payload53;
output 	src_payload54;
output 	src_payload55;
output 	src_payload56;
output 	src_payload57;
output 	src_payload58;
output 	src_payload59;
input 	last_write_collision;
input 	last_write_data_0;
input 	control_2;
input 	control_0;
output 	ShiftLeft1;
input 	last_write_data_1;
output 	ShiftLeft11;
input 	last_write_data_2;
output 	ShiftLeft12;
input 	last_write_data_3;
output 	ShiftLeft13;
input 	last_write_data_4;
output 	ShiftLeft14;
input 	last_write_data_5;
output 	ShiftLeft15;
input 	last_write_data_6;
output 	ShiftLeft16;
input 	last_write_data_7;
output 	ShiftLeft17;
input 	write_writedata;
input 	last_write_data_8;
output 	ShiftLeft18;
input 	write_writedata1;
input 	last_write_data_9;
output 	ShiftLeft19;
input 	write_writedata2;
input 	last_write_data_10;
output 	ShiftLeft110;
input 	write_writedata3;
input 	last_write_data_11;
output 	ShiftLeft111;
input 	write_writedata4;
input 	last_write_data_12;
output 	ShiftLeft112;
input 	write_writedata5;
input 	last_write_data_13;
output 	ShiftLeft113;
input 	write_writedata6;
input 	last_write_data_14;
output 	ShiftLeft114;
input 	write_writedata7;
input 	last_write_data_15;
output 	ShiftLeft115;
input 	last_write_data_16;
output 	ShiftLeft116;
input 	last_write_data_17;
output 	ShiftLeft117;
input 	last_write_data_18;
output 	ShiftLeft118;
input 	last_write_data_19;
output 	ShiftLeft119;
input 	last_write_data_20;
output 	ShiftLeft120;
input 	last_write_data_21;
output 	ShiftLeft121;
input 	last_write_data_22;
output 	ShiftLeft122;
input 	last_write_data_23;
output 	ShiftLeft123;
input 	last_write_data_24;
output 	ShiftLeft124;
input 	last_write_data_25;
output 	ShiftLeft125;
input 	last_write_data_26;
output 	ShiftLeft126;
input 	last_write_data_27;
output 	ShiftLeft127;
input 	last_write_data_28;
output 	ShiftLeft128;
input 	last_write_data_29;
output 	ShiftLeft129;
input 	last_write_data_30;
output 	ShiftLeft130;
input 	last_write_data_31;
output 	ShiftLeft131;
output 	ShiftLeft132;
output 	ShiftLeft133;
output 	ShiftLeft134;
output 	ShiftLeft135;
output 	ShiftLeft136;
output 	ShiftLeft137;
output 	ShiftLeft138;
output 	ShiftLeft139;
output 	ShiftLeft140;
output 	ShiftLeft141;
output 	ShiftLeft142;
output 	ShiftLeft143;
output 	ShiftLeft144;
output 	ShiftLeft145;
output 	ShiftLeft146;
output 	ShiftLeft147;
output 	ShiftLeft148;
output 	ShiftLeft149;
output 	ShiftLeft150;
output 	ShiftLeft151;
output 	ShiftLeft152;
output 	ShiftLeft153;
output 	ShiftLeft154;
output 	ShiftLeft155;
output 	ShiftLeft156;
output 	ShiftLeft157;
output 	ShiftLeft158;
output 	ShiftLeft159;
output 	ShiftLeft160;
output 	ShiftLeft161;
output 	ShiftLeft162;
output 	ShiftLeft163;
output 	ShiftLeft0;
output 	ShiftLeft01;
output 	ShiftLeft02;
output 	ShiftLeft03;
output 	ShiftLeft04;
output 	ShiftLeft05;
output 	ShiftLeft06;
output 	ShiftLeft07;
input 	altera_reset_synchronizer_int_chain_out;
output 	WideOr1;
input 	r_sync_rst;
input 	inc_read;
output 	av_readdatavalid;
output 	av_readdatavalid1;
output 	av_readdatavalid2;
output 	av_readdatavalid3;
input 	fifo_read;
output 	write_cp_ready;
output 	av_readdatavalid4;
output 	src0_valid;
output 	src_data_8;
output 	src_data_81;
output 	src_data_16;
output 	src_data_24;
output 	src_data_0;
output 	src_data_01;
output 	src_data_9;
output 	src_data_91;
output 	src_data_17;
output 	src_data_25;
output 	src_data_1;
output 	src_data_11;
output 	src_data_10;
output 	src_data_101;
output 	src_data_18;
output 	src_data_26;
output 	src_data_2;
output 	src_data_21;
output 	src_data_111;
output 	src_data_112;
output 	src_data_19;
output 	src_data_27;
output 	src_data_3;
output 	src_data_31;
output 	src_data_12;
output 	src_data_121;
output 	src_data_20;
output 	src_data_28;
output 	src_data_4;
output 	src_data_41;
output 	src_data_13;
output 	src_data_131;
output 	src_data_211;
output 	src_data_29;
output 	src_data_5;
output 	src_data_51;
output 	src_data_14;
output 	src_data_141;
output 	src_data_22;
output 	src_data_30;
output 	src_data_6;
output 	src_data_61;
output 	src_data_15;
output 	src_data_151;
output 	src_data_23;
output 	src_data_311;
output 	src_data_7;
output 	src_data_71;
output 	src_data_82;
output 	src_data_92;
output 	src_data_102;
output 	src_data_113;
output 	src_data_122;
output 	src_data_132;
output 	src_data_142;
output 	src_data_152;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][105]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][113]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][139]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][68]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][64]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][69]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][65]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][70]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][66]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][71]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][67]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][68]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][64]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][8]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][40]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][16]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][48]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][24]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][56]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][0]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][32]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][9]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][41]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][17]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][49]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][25]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][57]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][1]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][33]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][10]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][42]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][18]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][50]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][26]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][58]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][2]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][34]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][11]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][43]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][19]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][51]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][27]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][59]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][3]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][35]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][12]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][44]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][20]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][52]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][28]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][60]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][4]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][36]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][13]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][45]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][21]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][53]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][29]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][61]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][5]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][37]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][14]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][46]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][22]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][54]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][30]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][62]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][6]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][38]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][15]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][47]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][23]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][55]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][31]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][63]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][7]~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][39]~q ;
wire \dma_1_read_master_limiter|last_channel[1]~q ;
wire \dma_1_read_master_limiter|has_pending_responses~q ;
wire \arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[0]~q ;
wire \cmd_mux|src_payload~30_combout ;
wire \rsp_demux|src0_valid~0_combout ;
wire \arm_a9_hps_f2h_axi_slave_agent|bready~1_combout ;
wire \cmd_mux|src_payload~31_combout ;
wire \arm_a9_hps_f2h_axi_slave_rd_cmd_width_adapter|ShiftLeft0~0_combout ;


Computer_System_Computer_System_mm_interconnect_1_cmd_mux cmd_mux(
	.outclk_wire_0(outclk_wire_0),
	.writeaddress_2(writeaddress_2),
	.writeaddress_3(writeaddress_3),
	.writeaddress_4(writeaddress_4),
	.writeaddress_5(writeaddress_5),
	.writeaddress_6(writeaddress_6),
	.writeaddress_7(writeaddress_7),
	.writeaddress_8(writeaddress_8),
	.writeaddress_9(writeaddress_9),
	.writeaddress_10(writeaddress_10),
	.writeaddress_11(writeaddress_11),
	.writeaddress_12(writeaddress_12),
	.writeaddress_13(writeaddress_13),
	.writeaddress_14(writeaddress_14),
	.writeaddress_15(writeaddress_15),
	.writeaddress_16(writeaddress_16),
	.writeaddress_17(writeaddress_17),
	.writeaddress_18(writeaddress_18),
	.writeaddress_19(writeaddress_19),
	.writeaddress_20(writeaddress_20),
	.writeaddress_21(writeaddress_21),
	.writeaddress_22(writeaddress_22),
	.writeaddress_23(writeaddress_23),
	.writeaddress_24(writeaddress_24),
	.writeaddress_25(writeaddress_25),
	.writeaddress_26(writeaddress_26),
	.writeaddress_27(writeaddress_27),
	.writeaddress_28(writeaddress_28),
	.writeaddress_29(writeaddress_29),
	.writeaddress_30(writeaddress_30),
	.writeaddress_31(writeaddress_31),
	.hold_waitrequest(hold_waitrequest),
	.fifo_empty(fifo_empty),
	.saved_grant_1(saved_grant_1),
	.src_valid(src_valid),
	.src_payload(src_payload30),
	.src_payload1(src_payload31),
	.src_payload2(src_payload32),
	.src_payload3(src_payload33),
	.src_payload4(src_payload34),
	.src_payload5(src_payload35),
	.src_payload6(src_payload36),
	.src_payload7(src_payload37),
	.src_payload8(src_payload38),
	.src_payload9(src_payload39),
	.src_payload10(src_payload40),
	.src_payload11(src_payload41),
	.src_payload12(src_payload42),
	.src_payload13(src_payload43),
	.src_payload14(src_payload44),
	.src_payload15(src_payload45),
	.src_payload16(src_payload46),
	.src_payload17(src_payload47),
	.src_payload18(src_payload48),
	.src_payload19(src_payload49),
	.src_payload20(src_payload50),
	.src_payload21(src_payload51),
	.src_payload22(src_payload52),
	.src_payload23(src_payload53),
	.src_payload24(src_payload54),
	.src_payload25(src_payload55),
	.src_payload26(src_payload56),
	.src_payload27(src_payload57),
	.src_payload28(src_payload58),
	.src_payload29(src_payload59),
	.control_2(control_2),
	.control_0(control_0),
	.src_payload30(\cmd_mux|src_payload~30_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.write_cp_ready(write_cp_ready),
	.src_payload31(\cmd_mux|src_payload~31_combout ));

Computer_System_altera_merlin_traffic_limiter_2 dma_1_read_master_limiter(
	.f2h_BVALID_0(f2h_BVALID_0),
	.f2h_RVALID_0(f2h_RVALID_0),
	.clk(outclk_wire_0),
	.mem_105_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][105]~q ),
	.mem_113_0(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][113]~q ),
	.mem_139_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][139]~q ),
	.last_channel_1(\dma_1_read_master_limiter|last_channel[1]~q ),
	.has_pending_responses1(\dma_1_read_master_limiter|has_pending_responses~q ),
	.mem_used_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[0]~q ),
	.WideOr1(WideOr1),
	.reset(r_sync_rst),
	.inc_read(inc_read),
	.bready(\arm_a9_hps_f2h_axi_slave_agent|bready~1_combout ));

Computer_System_altera_merlin_axi_slave_ni arm_a9_hps_f2h_axi_slave_agent(
	.f2h_ARREADY_0(f2h_ARREADY_0),
	.f2h_AWREADY_0(f2h_AWREADY_0),
	.f2h_BVALID_0(f2h_BVALID_0),
	.f2h_RVALID_0(f2h_RVALID_0),
	.f2h_WREADY_0(f2h_WREADY_0),
	.outclk_wire_0(outclk_wire_0),
	.mem_105_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][105]~q ),
	.mem_113_0(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][113]~q ),
	.mem_139_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][139]~q ),
	.mem_68_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][68]~q ),
	.mem_64_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][64]~q ),
	.mem_69_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][69]~q ),
	.mem_65_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][65]~q ),
	.mem_70_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][70]~q ),
	.mem_66_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][66]~q ),
	.mem_71_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][71]~q ),
	.mem_67_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][67]~q ),
	.mem_68_01(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][68]~q ),
	.mem_64_01(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][64]~q ),
	.mem_8_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][8]~q ),
	.mem_40_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][40]~q ),
	.mem_16_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][16]~q ),
	.mem_48_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][48]~q ),
	.mem_24_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][24]~q ),
	.mem_56_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][56]~q ),
	.mem_0_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][0]~q ),
	.mem_32_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][32]~q ),
	.mem_9_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][9]~q ),
	.mem_41_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][41]~q ),
	.mem_17_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][17]~q ),
	.mem_49_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][49]~q ),
	.mem_25_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][25]~q ),
	.mem_57_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][57]~q ),
	.mem_1_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][1]~q ),
	.mem_33_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][33]~q ),
	.mem_10_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][10]~q ),
	.mem_42_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][42]~q ),
	.mem_18_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][18]~q ),
	.mem_50_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][50]~q ),
	.mem_26_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][26]~q ),
	.mem_58_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][58]~q ),
	.mem_2_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][2]~q ),
	.mem_34_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][34]~q ),
	.mem_11_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][11]~q ),
	.mem_43_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][43]~q ),
	.mem_19_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][19]~q ),
	.mem_51_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][51]~q ),
	.mem_27_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][27]~q ),
	.mem_59_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][59]~q ),
	.mem_3_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][3]~q ),
	.mem_35_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][35]~q ),
	.mem_12_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][12]~q ),
	.mem_44_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][44]~q ),
	.mem_20_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][20]~q ),
	.mem_52_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][52]~q ),
	.mem_28_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][28]~q ),
	.mem_60_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][60]~q ),
	.mem_4_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][4]~q ),
	.mem_36_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][36]~q ),
	.mem_13_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][13]~q ),
	.mem_45_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][45]~q ),
	.mem_21_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][21]~q ),
	.mem_53_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][53]~q ),
	.mem_29_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][29]~q ),
	.mem_61_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][61]~q ),
	.mem_5_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][5]~q ),
	.mem_37_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][37]~q ),
	.mem_14_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][14]~q ),
	.mem_46_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][46]~q ),
	.mem_22_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][22]~q ),
	.mem_54_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][54]~q ),
	.mem_30_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][30]~q ),
	.mem_62_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][62]~q ),
	.mem_6_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][6]~q ),
	.mem_38_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][38]~q ),
	.mem_15_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][15]~q ),
	.mem_47_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][47]~q ),
	.mem_23_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][23]~q ),
	.mem_55_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][55]~q ),
	.mem_31_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][31]~q ),
	.mem_63_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][63]~q ),
	.mem_7_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][7]~q ),
	.mem_39_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][39]~q ),
	.mem_used_7(mem_used_7),
	.saved_grant_0(saved_grant_0),
	.last_channel_1(\dma_1_read_master_limiter|last_channel[1]~q ),
	.has_pending_responses(\dma_1_read_master_limiter|has_pending_responses~q ),
	.read_select(read_select),
	.hold_waitrequest(hold_waitrequest),
	.write(write),
	.arvalid1(arvalid),
	.address_taken1(address_taken),
	.mem_used_71(mem_used_71),
	.saved_grant_1(saved_grant_1),
	.src_valid(src_valid),
	.awvalid1(awvalid),
	.mem_used_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[0]~q ),
	.bready(ARM_A9_HPS_f2h_axi_slave_bready),
	.data_taken1(data_taken),
	.wvalid1(wvalid),
	.src_payload(src_payload),
	.ShiftLeft1(ShiftLeft1),
	.ShiftLeft11(ShiftLeft11),
	.ShiftLeft12(ShiftLeft12),
	.ShiftLeft13(ShiftLeft13),
	.ShiftLeft14(ShiftLeft14),
	.ShiftLeft15(ShiftLeft15),
	.ShiftLeft16(ShiftLeft16),
	.ShiftLeft17(ShiftLeft17),
	.ShiftLeft18(ShiftLeft18),
	.ShiftLeft19(ShiftLeft19),
	.ShiftLeft110(ShiftLeft110),
	.ShiftLeft111(ShiftLeft111),
	.ShiftLeft112(ShiftLeft112),
	.ShiftLeft113(ShiftLeft113),
	.ShiftLeft114(ShiftLeft114),
	.ShiftLeft115(ShiftLeft115),
	.ShiftLeft116(ShiftLeft116),
	.ShiftLeft117(ShiftLeft117),
	.ShiftLeft118(ShiftLeft118),
	.ShiftLeft119(ShiftLeft119),
	.ShiftLeft120(ShiftLeft120),
	.ShiftLeft121(ShiftLeft121),
	.ShiftLeft122(ShiftLeft122),
	.ShiftLeft123(ShiftLeft123),
	.ShiftLeft124(ShiftLeft124),
	.ShiftLeft125(ShiftLeft125),
	.ShiftLeft126(ShiftLeft126),
	.ShiftLeft127(ShiftLeft127),
	.ShiftLeft128(ShiftLeft128),
	.ShiftLeft129(ShiftLeft129),
	.ShiftLeft130(ShiftLeft130),
	.ShiftLeft131(ShiftLeft131),
	.ShiftLeft132(ShiftLeft132),
	.ShiftLeft133(ShiftLeft133),
	.ShiftLeft134(ShiftLeft134),
	.ShiftLeft135(ShiftLeft135),
	.ShiftLeft136(ShiftLeft136),
	.ShiftLeft137(ShiftLeft137),
	.ShiftLeft138(ShiftLeft138),
	.ShiftLeft139(ShiftLeft139),
	.ShiftLeft140(ShiftLeft140),
	.ShiftLeft141(ShiftLeft141),
	.ShiftLeft142(ShiftLeft142),
	.ShiftLeft143(ShiftLeft143),
	.ShiftLeft144(ShiftLeft144),
	.ShiftLeft145(ShiftLeft145),
	.ShiftLeft146(ShiftLeft146),
	.ShiftLeft147(ShiftLeft147),
	.ShiftLeft148(ShiftLeft148),
	.ShiftLeft149(ShiftLeft149),
	.ShiftLeft150(ShiftLeft150),
	.ShiftLeft151(ShiftLeft151),
	.ShiftLeft152(ShiftLeft152),
	.ShiftLeft153(ShiftLeft153),
	.ShiftLeft154(ShiftLeft154),
	.ShiftLeft155(ShiftLeft155),
	.ShiftLeft156(ShiftLeft156),
	.ShiftLeft157(ShiftLeft157),
	.ShiftLeft158(ShiftLeft158),
	.ShiftLeft159(ShiftLeft159),
	.ShiftLeft160(ShiftLeft160),
	.ShiftLeft161(ShiftLeft161),
	.ShiftLeft162(ShiftLeft162),
	.ShiftLeft163(ShiftLeft163),
	.ShiftLeft0(ShiftLeft0),
	.ShiftLeft01(ShiftLeft01),
	.ShiftLeft02(ShiftLeft02),
	.ShiftLeft03(ShiftLeft03),
	.ShiftLeft04(ShiftLeft04),
	.ShiftLeft05(ShiftLeft05),
	.ShiftLeft06(ShiftLeft06),
	.ShiftLeft07(ShiftLeft07),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.fifo_read(fifo_read),
	.bready1(\arm_a9_hps_f2h_axi_slave_agent|bready~1_combout ),
	.write_cp_ready(write_cp_ready),
	.src_payload1(\cmd_mux|src_payload~31_combout ),
	.ShiftLeft08(\arm_a9_hps_f2h_axi_slave_rd_cmd_width_adapter|ShiftLeft0~0_combout ));

Computer_System_altera_merlin_master_agent dma_1_read_master_agent(
	.f2h_BVALID_0(f2h_BVALID_0),
	.f2h_RVALID_0(f2h_RVALID_0),
	.mem_68_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][68]~q ),
	.mem_64_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][64]~q ),
	.mem_69_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][69]~q ),
	.mem_65_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][65]~q ),
	.mem_70_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][70]~q ),
	.mem_66_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][66]~q ),
	.mem_71_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][71]~q ),
	.mem_67_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][67]~q ),
	.mem_68_01(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][68]~q ),
	.mem_64_01(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][64]~q ),
	.mem_used_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[0]~q ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.av_readdatavalid(av_readdatavalid),
	.av_readdatavalid1(av_readdatavalid1),
	.av_readdatavalid2(av_readdatavalid2),
	.av_readdatavalid3(av_readdatavalid3),
	.av_readdatavalid4(av_readdatavalid4));

Computer_System_Computer_System_mm_interconnect_1_rsp_mux rsp_mux(
	.f2h_BVALID_0(f2h_BVALID_0),
	.f2h_RVALID_0(f2h_RVALID_0),
	.f2h_RDATA_0(f2h_RDATA_0),
	.f2h_RDATA_1(f2h_RDATA_1),
	.f2h_RDATA_2(f2h_RDATA_2),
	.f2h_RDATA_3(f2h_RDATA_3),
	.f2h_RDATA_4(f2h_RDATA_4),
	.f2h_RDATA_5(f2h_RDATA_5),
	.f2h_RDATA_6(f2h_RDATA_6),
	.f2h_RDATA_7(f2h_RDATA_7),
	.f2h_RDATA_8(f2h_RDATA_8),
	.f2h_RDATA_9(f2h_RDATA_9),
	.f2h_RDATA_10(f2h_RDATA_10),
	.f2h_RDATA_11(f2h_RDATA_11),
	.f2h_RDATA_12(f2h_RDATA_12),
	.f2h_RDATA_13(f2h_RDATA_13),
	.f2h_RDATA_14(f2h_RDATA_14),
	.f2h_RDATA_15(f2h_RDATA_15),
	.f2h_RDATA_16(f2h_RDATA_16),
	.f2h_RDATA_17(f2h_RDATA_17),
	.f2h_RDATA_18(f2h_RDATA_18),
	.f2h_RDATA_19(f2h_RDATA_19),
	.f2h_RDATA_20(f2h_RDATA_20),
	.f2h_RDATA_21(f2h_RDATA_21),
	.f2h_RDATA_22(f2h_RDATA_22),
	.f2h_RDATA_23(f2h_RDATA_23),
	.f2h_RDATA_24(f2h_RDATA_24),
	.f2h_RDATA_25(f2h_RDATA_25),
	.f2h_RDATA_26(f2h_RDATA_26),
	.f2h_RDATA_27(f2h_RDATA_27),
	.f2h_RDATA_28(f2h_RDATA_28),
	.f2h_RDATA_29(f2h_RDATA_29),
	.f2h_RDATA_30(f2h_RDATA_30),
	.f2h_RDATA_31(f2h_RDATA_31),
	.f2h_RDATA_32(f2h_RDATA_32),
	.f2h_RDATA_33(f2h_RDATA_33),
	.f2h_RDATA_34(f2h_RDATA_34),
	.f2h_RDATA_35(f2h_RDATA_35),
	.f2h_RDATA_36(f2h_RDATA_36),
	.f2h_RDATA_37(f2h_RDATA_37),
	.f2h_RDATA_38(f2h_RDATA_38),
	.f2h_RDATA_39(f2h_RDATA_39),
	.f2h_RDATA_40(f2h_RDATA_40),
	.f2h_RDATA_41(f2h_RDATA_41),
	.f2h_RDATA_42(f2h_RDATA_42),
	.f2h_RDATA_43(f2h_RDATA_43),
	.f2h_RDATA_44(f2h_RDATA_44),
	.f2h_RDATA_45(f2h_RDATA_45),
	.f2h_RDATA_46(f2h_RDATA_46),
	.f2h_RDATA_47(f2h_RDATA_47),
	.f2h_RDATA_48(f2h_RDATA_48),
	.f2h_RDATA_49(f2h_RDATA_49),
	.f2h_RDATA_50(f2h_RDATA_50),
	.f2h_RDATA_51(f2h_RDATA_51),
	.f2h_RDATA_52(f2h_RDATA_52),
	.f2h_RDATA_53(f2h_RDATA_53),
	.f2h_RDATA_54(f2h_RDATA_54),
	.f2h_RDATA_55(f2h_RDATA_55),
	.f2h_RDATA_56(f2h_RDATA_56),
	.f2h_RDATA_57(f2h_RDATA_57),
	.f2h_RDATA_58(f2h_RDATA_58),
	.f2h_RDATA_59(f2h_RDATA_59),
	.f2h_RDATA_60(f2h_RDATA_60),
	.f2h_RDATA_61(f2h_RDATA_61),
	.f2h_RDATA_62(f2h_RDATA_62),
	.f2h_RDATA_63(f2h_RDATA_63),
	.mem_68_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][68]~q ),
	.mem_64_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][64]~q ),
	.mem_69_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][69]~q ),
	.mem_65_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][65]~q ),
	.mem_70_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][70]~q ),
	.mem_66_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][66]~q ),
	.mem_71_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][71]~q ),
	.mem_67_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][67]~q ),
	.mem_68_01(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][68]~q ),
	.mem_64_01(\arm_a9_hps_f2h_axi_slave_agent|read_rsp_fifo|mem[0][64]~q ),
	.mem_8_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][8]~q ),
	.mem_40_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][40]~q ),
	.mem_16_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][16]~q ),
	.mem_48_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][48]~q ),
	.mem_24_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][24]~q ),
	.mem_56_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][56]~q ),
	.mem_0_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][0]~q ),
	.mem_32_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][32]~q ),
	.mem_9_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][9]~q ),
	.mem_41_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][41]~q ),
	.mem_17_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][17]~q ),
	.mem_49_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][49]~q ),
	.mem_25_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][25]~q ),
	.mem_57_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][57]~q ),
	.mem_1_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][1]~q ),
	.mem_33_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][33]~q ),
	.mem_10_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][10]~q ),
	.mem_42_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][42]~q ),
	.mem_18_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][18]~q ),
	.mem_50_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][50]~q ),
	.mem_26_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][26]~q ),
	.mem_58_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][58]~q ),
	.mem_2_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][2]~q ),
	.mem_34_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][34]~q ),
	.mem_11_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][11]~q ),
	.mem_43_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][43]~q ),
	.mem_19_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][19]~q ),
	.mem_51_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][51]~q ),
	.mem_27_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][27]~q ),
	.mem_59_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][59]~q ),
	.mem_3_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][3]~q ),
	.mem_35_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][35]~q ),
	.mem_12_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][12]~q ),
	.mem_44_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][44]~q ),
	.mem_20_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][20]~q ),
	.mem_52_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][52]~q ),
	.mem_28_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][28]~q ),
	.mem_60_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][60]~q ),
	.mem_4_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][4]~q ),
	.mem_36_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][36]~q ),
	.mem_13_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][13]~q ),
	.mem_45_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][45]~q ),
	.mem_21_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][21]~q ),
	.mem_53_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][53]~q ),
	.mem_29_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][29]~q ),
	.mem_61_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][61]~q ),
	.mem_5_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][5]~q ),
	.mem_37_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][37]~q ),
	.mem_14_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][14]~q ),
	.mem_46_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][46]~q ),
	.mem_22_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][22]~q ),
	.mem_54_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][54]~q ),
	.mem_30_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][30]~q ),
	.mem_62_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][62]~q ),
	.mem_6_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][6]~q ),
	.mem_38_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][38]~q ),
	.mem_15_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][15]~q ),
	.mem_47_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][47]~q ),
	.mem_23_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][23]~q ),
	.mem_55_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][55]~q ),
	.mem_31_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][31]~q ),
	.mem_63_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][63]~q ),
	.mem_7_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][7]~q ),
	.mem_39_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][39]~q ),
	.mem_used_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[0]~q ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.src_data_8(src_data_8),
	.src_data_81(src_data_81),
	.src_data_16(src_data_16),
	.src_data_24(src_data_24),
	.src_data_0(src_data_0),
	.src_data_01(src_data_01),
	.src_data_9(src_data_9),
	.src_data_91(src_data_91),
	.src_data_17(src_data_17),
	.src_data_25(src_data_25),
	.src_data_1(src_data_1),
	.src_data_11(src_data_11),
	.src_data_10(src_data_10),
	.src_data_101(src_data_101),
	.src_data_18(src_data_18),
	.src_data_26(src_data_26),
	.src_data_2(src_data_2),
	.src_data_21(src_data_21),
	.src_data_111(src_data_111),
	.src_data_112(src_data_112),
	.src_data_19(src_data_19),
	.src_data_27(src_data_27),
	.src_data_3(src_data_3),
	.src_data_31(src_data_31),
	.src_data_12(src_data_12),
	.src_data_121(src_data_121),
	.src_data_20(src_data_20),
	.src_data_28(src_data_28),
	.src_data_4(src_data_4),
	.src_data_41(src_data_41),
	.src_data_13(src_data_13),
	.src_data_131(src_data_131),
	.src_data_211(src_data_211),
	.src_data_29(src_data_29),
	.src_data_5(src_data_5),
	.src_data_51(src_data_51),
	.src_data_14(src_data_14),
	.src_data_141(src_data_141),
	.src_data_22(src_data_22),
	.src_data_30(src_data_30),
	.src_data_6(src_data_6),
	.src_data_61(src_data_61),
	.src_data_15(src_data_15),
	.src_data_151(src_data_151),
	.src_data_23(src_data_23),
	.src_data_311(src_data_311),
	.src_data_7(src_data_7),
	.src_data_71(src_data_71),
	.src_data_82(src_data_82),
	.src_data_92(src_data_92),
	.src_data_102(src_data_102),
	.src_data_113(src_data_113),
	.src_data_122(src_data_122),
	.src_data_132(src_data_132),
	.src_data_142(src_data_142),
	.src_data_152(src_data_152));

Computer_System_Computer_System_mm_interconnect_1_cmd_demux_001_1 rsp_demux(
	.f2h_BVALID_0(f2h_BVALID_0),
	.mem_105_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][105]~q ),
	.mem_139_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem[0][139]~q ),
	.mem_used_0(\arm_a9_hps_f2h_axi_slave_agent|write_rsp_fifo|mem_used[0]~q ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.src0_valid1(src0_valid));

Computer_System_Computer_System_mm_interconnect_1_cmd_mux_1 cmd_mux_001(
	.f2h_ARREADY_0(f2h_ARREADY_0),
	.outclk_wire_0(outclk_wire_0),
	.readaddress_2(readaddress_2),
	.readaddress_3(readaddress_3),
	.readaddress_4(readaddress_4),
	.readaddress_5(readaddress_5),
	.readaddress_6(readaddress_6),
	.readaddress_7(readaddress_7),
	.readaddress_8(readaddress_8),
	.readaddress_9(readaddress_9),
	.readaddress_10(readaddress_10),
	.readaddress_11(readaddress_11),
	.readaddress_12(readaddress_12),
	.readaddress_13(readaddress_13),
	.readaddress_14(readaddress_14),
	.readaddress_15(readaddress_15),
	.readaddress_16(readaddress_16),
	.readaddress_17(readaddress_17),
	.readaddress_18(readaddress_18),
	.readaddress_19(readaddress_19),
	.readaddress_20(readaddress_20),
	.readaddress_21(readaddress_21),
	.readaddress_22(readaddress_22),
	.readaddress_23(readaddress_23),
	.readaddress_24(readaddress_24),
	.readaddress_25(readaddress_25),
	.readaddress_26(readaddress_26),
	.readaddress_27(readaddress_27),
	.readaddress_28(readaddress_28),
	.readaddress_29(readaddress_29),
	.readaddress_30(readaddress_30),
	.readaddress_31(readaddress_31),
	.mem_used_7(mem_used_7),
	.saved_grant_0(saved_grant_0),
	.last_channel_1(\dma_1_read_master_limiter|last_channel[1]~q ),
	.has_pending_responses(\dma_1_read_master_limiter|has_pending_responses~q ),
	.read_select(read_select),
	.hold_waitrequest(hold_waitrequest),
	.write(write),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.WideOr1(WideOr1));

Computer_System_altera_merlin_width_adapter arm_a9_hps_f2h_axi_slave_rd_cmd_width_adapter(
	.readaddress_2(readaddress_2),
	.saved_grant_0(saved_grant_0),
	.ShiftLeft0(\arm_a9_hps_f2h_axi_slave_rd_cmd_width_adapter|ShiftLeft0~0_combout ));

Computer_System_altera_merlin_width_adapter_2 arm_a9_hps_f2h_axi_slave_wr_cmd_width_adapter(
	.writeaddress_2(writeaddress_2),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.writeaddress_1(writeaddress_1),
	.writeaddress_0(writeaddress_0),
	.saved_grant_1(saved_grant_1),
	.last_write_collision(last_write_collision),
	.last_write_data_0(last_write_data_0),
	.control_2(control_2),
	.control_0(control_0),
	.src_payload(\cmd_mux|src_payload~30_combout ),
	.ShiftLeft1(ShiftLeft1),
	.last_write_data_1(last_write_data_1),
	.ShiftLeft11(ShiftLeft11),
	.last_write_data_2(last_write_data_2),
	.ShiftLeft12(ShiftLeft12),
	.last_write_data_3(last_write_data_3),
	.ShiftLeft13(ShiftLeft13),
	.last_write_data_4(last_write_data_4),
	.ShiftLeft14(ShiftLeft14),
	.last_write_data_5(last_write_data_5),
	.ShiftLeft15(ShiftLeft15),
	.last_write_data_6(last_write_data_6),
	.ShiftLeft16(ShiftLeft16),
	.last_write_data_7(last_write_data_7),
	.ShiftLeft17(ShiftLeft17),
	.write_writedata(write_writedata),
	.last_write_data_8(last_write_data_8),
	.ShiftLeft18(ShiftLeft18),
	.write_writedata1(write_writedata1),
	.last_write_data_9(last_write_data_9),
	.ShiftLeft19(ShiftLeft19),
	.write_writedata2(write_writedata2),
	.last_write_data_10(last_write_data_10),
	.ShiftLeft110(ShiftLeft110),
	.write_writedata3(write_writedata3),
	.last_write_data_11(last_write_data_11),
	.ShiftLeft111(ShiftLeft111),
	.write_writedata4(write_writedata4),
	.last_write_data_12(last_write_data_12),
	.ShiftLeft112(ShiftLeft112),
	.write_writedata5(write_writedata5),
	.last_write_data_13(last_write_data_13),
	.ShiftLeft113(ShiftLeft113),
	.write_writedata6(write_writedata6),
	.last_write_data_14(last_write_data_14),
	.ShiftLeft114(ShiftLeft114),
	.write_writedata7(write_writedata7),
	.last_write_data_15(last_write_data_15),
	.ShiftLeft115(ShiftLeft115),
	.last_write_data_16(last_write_data_16),
	.ShiftLeft116(ShiftLeft116),
	.last_write_data_17(last_write_data_17),
	.ShiftLeft117(ShiftLeft117),
	.last_write_data_18(last_write_data_18),
	.ShiftLeft118(ShiftLeft118),
	.last_write_data_19(last_write_data_19),
	.ShiftLeft119(ShiftLeft119),
	.last_write_data_20(last_write_data_20),
	.ShiftLeft120(ShiftLeft120),
	.last_write_data_21(last_write_data_21),
	.ShiftLeft121(ShiftLeft121),
	.last_write_data_22(last_write_data_22),
	.ShiftLeft122(ShiftLeft122),
	.last_write_data_23(last_write_data_23),
	.ShiftLeft123(ShiftLeft123),
	.last_write_data_24(last_write_data_24),
	.ShiftLeft124(ShiftLeft124),
	.last_write_data_25(last_write_data_25),
	.ShiftLeft125(ShiftLeft125),
	.last_write_data_26(last_write_data_26),
	.ShiftLeft126(ShiftLeft126),
	.last_write_data_27(last_write_data_27),
	.ShiftLeft127(ShiftLeft127),
	.last_write_data_28(last_write_data_28),
	.ShiftLeft128(ShiftLeft128),
	.last_write_data_29(last_write_data_29),
	.ShiftLeft129(ShiftLeft129),
	.last_write_data_30(last_write_data_30),
	.ShiftLeft130(ShiftLeft130),
	.last_write_data_31(last_write_data_31),
	.ShiftLeft131(ShiftLeft131),
	.ShiftLeft132(ShiftLeft132),
	.ShiftLeft133(ShiftLeft133),
	.ShiftLeft134(ShiftLeft134),
	.ShiftLeft135(ShiftLeft135),
	.ShiftLeft136(ShiftLeft136),
	.ShiftLeft137(ShiftLeft137),
	.ShiftLeft138(ShiftLeft138),
	.ShiftLeft139(ShiftLeft139),
	.ShiftLeft140(ShiftLeft140),
	.ShiftLeft141(ShiftLeft141),
	.ShiftLeft142(ShiftLeft142),
	.ShiftLeft143(ShiftLeft143),
	.ShiftLeft144(ShiftLeft144),
	.ShiftLeft145(ShiftLeft145),
	.ShiftLeft146(ShiftLeft146),
	.ShiftLeft147(ShiftLeft147),
	.ShiftLeft148(ShiftLeft148),
	.ShiftLeft149(ShiftLeft149),
	.ShiftLeft150(ShiftLeft150),
	.ShiftLeft151(ShiftLeft151),
	.ShiftLeft152(ShiftLeft152),
	.ShiftLeft153(ShiftLeft153),
	.ShiftLeft154(ShiftLeft154),
	.ShiftLeft155(ShiftLeft155),
	.ShiftLeft156(ShiftLeft156),
	.ShiftLeft157(ShiftLeft157),
	.ShiftLeft158(ShiftLeft158),
	.ShiftLeft159(ShiftLeft159),
	.ShiftLeft160(ShiftLeft160),
	.ShiftLeft161(ShiftLeft161),
	.ShiftLeft162(ShiftLeft162),
	.ShiftLeft163(ShiftLeft163),
	.ShiftLeft0(ShiftLeft0),
	.ShiftLeft01(ShiftLeft01),
	.ShiftLeft02(ShiftLeft02),
	.ShiftLeft03(ShiftLeft03),
	.ShiftLeft04(ShiftLeft04),
	.ShiftLeft05(ShiftLeft05),
	.ShiftLeft06(ShiftLeft06),
	.ShiftLeft07(ShiftLeft07));

endmodule

module Computer_System_altera_merlin_axi_slave_ni (
	f2h_ARREADY_0,
	f2h_AWREADY_0,
	f2h_BVALID_0,
	f2h_RVALID_0,
	f2h_WREADY_0,
	outclk_wire_0,
	mem_105_0,
	mem_113_0,
	mem_139_0,
	mem_68_0,
	mem_64_0,
	mem_69_0,
	mem_65_0,
	mem_70_0,
	mem_66_0,
	mem_71_0,
	mem_67_0,
	mem_68_01,
	mem_64_01,
	mem_8_0,
	mem_40_0,
	mem_16_0,
	mem_48_0,
	mem_24_0,
	mem_56_0,
	mem_0_0,
	mem_32_0,
	mem_9_0,
	mem_41_0,
	mem_17_0,
	mem_49_0,
	mem_25_0,
	mem_57_0,
	mem_1_0,
	mem_33_0,
	mem_10_0,
	mem_42_0,
	mem_18_0,
	mem_50_0,
	mem_26_0,
	mem_58_0,
	mem_2_0,
	mem_34_0,
	mem_11_0,
	mem_43_0,
	mem_19_0,
	mem_51_0,
	mem_27_0,
	mem_59_0,
	mem_3_0,
	mem_35_0,
	mem_12_0,
	mem_44_0,
	mem_20_0,
	mem_52_0,
	mem_28_0,
	mem_60_0,
	mem_4_0,
	mem_36_0,
	mem_13_0,
	mem_45_0,
	mem_21_0,
	mem_53_0,
	mem_29_0,
	mem_61_0,
	mem_5_0,
	mem_37_0,
	mem_14_0,
	mem_46_0,
	mem_22_0,
	mem_54_0,
	mem_30_0,
	mem_62_0,
	mem_6_0,
	mem_38_0,
	mem_15_0,
	mem_47_0,
	mem_23_0,
	mem_55_0,
	mem_31_0,
	mem_63_0,
	mem_7_0,
	mem_39_0,
	mem_used_7,
	saved_grant_0,
	last_channel_1,
	has_pending_responses,
	read_select,
	hold_waitrequest,
	write,
	arvalid1,
	address_taken1,
	mem_used_71,
	saved_grant_1,
	src_valid,
	awvalid1,
	mem_used_0,
	bready,
	data_taken1,
	wvalid1,
	src_payload,
	ShiftLeft1,
	ShiftLeft11,
	ShiftLeft12,
	ShiftLeft13,
	ShiftLeft14,
	ShiftLeft15,
	ShiftLeft16,
	ShiftLeft17,
	ShiftLeft18,
	ShiftLeft19,
	ShiftLeft110,
	ShiftLeft111,
	ShiftLeft112,
	ShiftLeft113,
	ShiftLeft114,
	ShiftLeft115,
	ShiftLeft116,
	ShiftLeft117,
	ShiftLeft118,
	ShiftLeft119,
	ShiftLeft120,
	ShiftLeft121,
	ShiftLeft122,
	ShiftLeft123,
	ShiftLeft124,
	ShiftLeft125,
	ShiftLeft126,
	ShiftLeft127,
	ShiftLeft128,
	ShiftLeft129,
	ShiftLeft130,
	ShiftLeft131,
	ShiftLeft132,
	ShiftLeft133,
	ShiftLeft134,
	ShiftLeft135,
	ShiftLeft136,
	ShiftLeft137,
	ShiftLeft138,
	ShiftLeft139,
	ShiftLeft140,
	ShiftLeft141,
	ShiftLeft142,
	ShiftLeft143,
	ShiftLeft144,
	ShiftLeft145,
	ShiftLeft146,
	ShiftLeft147,
	ShiftLeft148,
	ShiftLeft149,
	ShiftLeft150,
	ShiftLeft151,
	ShiftLeft152,
	ShiftLeft153,
	ShiftLeft154,
	ShiftLeft155,
	ShiftLeft156,
	ShiftLeft157,
	ShiftLeft158,
	ShiftLeft159,
	ShiftLeft160,
	ShiftLeft161,
	ShiftLeft162,
	ShiftLeft163,
	ShiftLeft0,
	ShiftLeft01,
	ShiftLeft02,
	ShiftLeft03,
	ShiftLeft04,
	ShiftLeft05,
	ShiftLeft06,
	ShiftLeft07,
	altera_reset_synchronizer_int_chain_out,
	fifo_read,
	bready1,
	write_cp_ready,
	src_payload1,
	ShiftLeft08)/* synthesis synthesis_greybox=0 */;
input 	f2h_ARREADY_0;
input 	f2h_AWREADY_0;
input 	f2h_BVALID_0;
input 	f2h_RVALID_0;
input 	f2h_WREADY_0;
input 	outclk_wire_0;
output 	mem_105_0;
output 	mem_113_0;
output 	mem_139_0;
output 	mem_68_0;
output 	mem_64_0;
output 	mem_69_0;
output 	mem_65_0;
output 	mem_70_0;
output 	mem_66_0;
output 	mem_71_0;
output 	mem_67_0;
output 	mem_68_01;
output 	mem_64_01;
output 	mem_8_0;
output 	mem_40_0;
output 	mem_16_0;
output 	mem_48_0;
output 	mem_24_0;
output 	mem_56_0;
output 	mem_0_0;
output 	mem_32_0;
output 	mem_9_0;
output 	mem_41_0;
output 	mem_17_0;
output 	mem_49_0;
output 	mem_25_0;
output 	mem_57_0;
output 	mem_1_0;
output 	mem_33_0;
output 	mem_10_0;
output 	mem_42_0;
output 	mem_18_0;
output 	mem_50_0;
output 	mem_26_0;
output 	mem_58_0;
output 	mem_2_0;
output 	mem_34_0;
output 	mem_11_0;
output 	mem_43_0;
output 	mem_19_0;
output 	mem_51_0;
output 	mem_27_0;
output 	mem_59_0;
output 	mem_3_0;
output 	mem_35_0;
output 	mem_12_0;
output 	mem_44_0;
output 	mem_20_0;
output 	mem_52_0;
output 	mem_28_0;
output 	mem_60_0;
output 	mem_4_0;
output 	mem_36_0;
output 	mem_13_0;
output 	mem_45_0;
output 	mem_21_0;
output 	mem_53_0;
output 	mem_29_0;
output 	mem_61_0;
output 	mem_5_0;
output 	mem_37_0;
output 	mem_14_0;
output 	mem_46_0;
output 	mem_22_0;
output 	mem_54_0;
output 	mem_30_0;
output 	mem_62_0;
output 	mem_6_0;
output 	mem_38_0;
output 	mem_15_0;
output 	mem_47_0;
output 	mem_23_0;
output 	mem_55_0;
output 	mem_31_0;
output 	mem_63_0;
output 	mem_7_0;
output 	mem_39_0;
output 	mem_used_7;
input 	saved_grant_0;
input 	last_channel_1;
input 	has_pending_responses;
input 	read_select;
input 	hold_waitrequest;
output 	write;
output 	arvalid1;
output 	address_taken1;
output 	mem_used_71;
input 	saved_grant_1;
input 	src_valid;
output 	awvalid1;
output 	mem_used_0;
output 	bready;
output 	data_taken1;
output 	wvalid1;
input 	src_payload;
input 	ShiftLeft1;
input 	ShiftLeft11;
input 	ShiftLeft12;
input 	ShiftLeft13;
input 	ShiftLeft14;
input 	ShiftLeft15;
input 	ShiftLeft16;
input 	ShiftLeft17;
input 	ShiftLeft18;
input 	ShiftLeft19;
input 	ShiftLeft110;
input 	ShiftLeft111;
input 	ShiftLeft112;
input 	ShiftLeft113;
input 	ShiftLeft114;
input 	ShiftLeft115;
input 	ShiftLeft116;
input 	ShiftLeft117;
input 	ShiftLeft118;
input 	ShiftLeft119;
input 	ShiftLeft120;
input 	ShiftLeft121;
input 	ShiftLeft122;
input 	ShiftLeft123;
input 	ShiftLeft124;
input 	ShiftLeft125;
input 	ShiftLeft126;
input 	ShiftLeft127;
input 	ShiftLeft128;
input 	ShiftLeft129;
input 	ShiftLeft130;
input 	ShiftLeft131;
input 	ShiftLeft132;
input 	ShiftLeft133;
input 	ShiftLeft134;
input 	ShiftLeft135;
input 	ShiftLeft136;
input 	ShiftLeft137;
input 	ShiftLeft138;
input 	ShiftLeft139;
input 	ShiftLeft140;
input 	ShiftLeft141;
input 	ShiftLeft142;
input 	ShiftLeft143;
input 	ShiftLeft144;
input 	ShiftLeft145;
input 	ShiftLeft146;
input 	ShiftLeft147;
input 	ShiftLeft148;
input 	ShiftLeft149;
input 	ShiftLeft150;
input 	ShiftLeft151;
input 	ShiftLeft152;
input 	ShiftLeft153;
input 	ShiftLeft154;
input 	ShiftLeft155;
input 	ShiftLeft156;
input 	ShiftLeft157;
input 	ShiftLeft158;
input 	ShiftLeft159;
input 	ShiftLeft160;
input 	ShiftLeft161;
input 	ShiftLeft162;
input 	ShiftLeft163;
input 	ShiftLeft0;
input 	ShiftLeft01;
input 	ShiftLeft02;
input 	ShiftLeft03;
input 	ShiftLeft04;
input 	ShiftLeft05;
input 	ShiftLeft06;
input 	ShiftLeft07;
input 	altera_reset_synchronizer_int_chain_out;
input 	fifo_read;
output 	bready1;
output 	write_cp_ready;
input 	src_payload1;
input 	ShiftLeft08;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_taken~0_combout ;
wire \data_taken~0_combout ;


Computer_System_altera_avalon_sc_fifo_4 read_rsp_fifo(
	.f2h_ARREADY_0(f2h_ARREADY_0),
	.f2h_RVALID_0(f2h_RVALID_0),
	.clk(outclk_wire_0),
	.mem_113_0(mem_113_0),
	.mem_68_0(mem_68_01),
	.mem_64_0(mem_64_01),
	.mem_used_7(mem_used_7),
	.saved_grant_0(saved_grant_0),
	.last_channel_1(last_channel_1),
	.has_pending_responses(has_pending_responses),
	.read_select(read_select),
	.hold_waitrequest(hold_waitrequest),
	.write(write),
	.src_payload(src_payload),
	.reset(altera_reset_synchronizer_int_chain_out),
	.ShiftLeft0(ShiftLeft08));

Computer_System_altera_avalon_sc_fifo_5 write_rsp_fifo(
	.f2h_BVALID_0(f2h_BVALID_0),
	.clk(outclk_wire_0),
	.mem_105_0(mem_105_0),
	.mem_139_0(mem_139_0),
	.mem_68_0(mem_68_0),
	.mem_64_0(mem_64_0),
	.mem_69_0(mem_69_0),
	.mem_65_0(mem_65_0),
	.mem_70_0(mem_70_0),
	.mem_66_0(mem_66_0),
	.mem_71_0(mem_71_0),
	.mem_67_0(mem_67_0),
	.mem_8_0(mem_8_0),
	.mem_40_0(mem_40_0),
	.mem_16_0(mem_16_0),
	.mem_48_0(mem_48_0),
	.mem_24_0(mem_24_0),
	.mem_56_0(mem_56_0),
	.mem_0_0(mem_0_0),
	.mem_32_0(mem_32_0),
	.mem_9_0(mem_9_0),
	.mem_41_0(mem_41_0),
	.mem_17_0(mem_17_0),
	.mem_49_0(mem_49_0),
	.mem_25_0(mem_25_0),
	.mem_57_0(mem_57_0),
	.mem_1_0(mem_1_0),
	.mem_33_0(mem_33_0),
	.mem_10_0(mem_10_0),
	.mem_42_0(mem_42_0),
	.mem_18_0(mem_18_0),
	.mem_50_0(mem_50_0),
	.mem_26_0(mem_26_0),
	.mem_58_0(mem_58_0),
	.mem_2_0(mem_2_0),
	.mem_34_0(mem_34_0),
	.mem_11_0(mem_11_0),
	.mem_43_0(mem_43_0),
	.mem_19_0(mem_19_0),
	.mem_51_0(mem_51_0),
	.mem_27_0(mem_27_0),
	.mem_59_0(mem_59_0),
	.mem_3_0(mem_3_0),
	.mem_35_0(mem_35_0),
	.mem_12_0(mem_12_0),
	.mem_44_0(mem_44_0),
	.mem_20_0(mem_20_0),
	.mem_52_0(mem_52_0),
	.mem_28_0(mem_28_0),
	.mem_60_0(mem_60_0),
	.mem_4_0(mem_4_0),
	.mem_36_0(mem_36_0),
	.mem_13_0(mem_13_0),
	.mem_45_0(mem_45_0),
	.mem_21_0(mem_21_0),
	.mem_53_0(mem_53_0),
	.mem_29_0(mem_29_0),
	.mem_61_0(mem_61_0),
	.mem_5_0(mem_5_0),
	.mem_37_0(mem_37_0),
	.mem_14_0(mem_14_0),
	.mem_46_0(mem_46_0),
	.mem_22_0(mem_22_0),
	.mem_54_0(mem_54_0),
	.mem_30_0(mem_30_0),
	.mem_62_0(mem_62_0),
	.mem_6_0(mem_6_0),
	.mem_38_0(mem_38_0),
	.mem_15_0(mem_15_0),
	.mem_47_0(mem_47_0),
	.mem_23_0(mem_23_0),
	.mem_55_0(mem_55_0),
	.mem_31_0(mem_31_0),
	.mem_63_0(mem_63_0),
	.mem_7_0(mem_7_0),
	.mem_39_0(mem_39_0),
	.mem_used_7(mem_used_71),
	.saved_grant_1(saved_grant_1),
	.src_valid(src_valid),
	.mem_used_0(mem_used_0),
	.ShiftLeft1(ShiftLeft1),
	.ShiftLeft11(ShiftLeft11),
	.ShiftLeft12(ShiftLeft12),
	.ShiftLeft13(ShiftLeft13),
	.ShiftLeft14(ShiftLeft14),
	.ShiftLeft15(ShiftLeft15),
	.ShiftLeft16(ShiftLeft16),
	.ShiftLeft17(ShiftLeft17),
	.ShiftLeft18(ShiftLeft18),
	.ShiftLeft19(ShiftLeft19),
	.ShiftLeft110(ShiftLeft110),
	.ShiftLeft111(ShiftLeft111),
	.ShiftLeft112(ShiftLeft112),
	.ShiftLeft113(ShiftLeft113),
	.ShiftLeft114(ShiftLeft114),
	.ShiftLeft115(ShiftLeft115),
	.ShiftLeft116(ShiftLeft116),
	.ShiftLeft117(ShiftLeft117),
	.ShiftLeft118(ShiftLeft118),
	.ShiftLeft119(ShiftLeft119),
	.ShiftLeft120(ShiftLeft120),
	.ShiftLeft121(ShiftLeft121),
	.ShiftLeft122(ShiftLeft122),
	.ShiftLeft123(ShiftLeft123),
	.ShiftLeft124(ShiftLeft124),
	.ShiftLeft125(ShiftLeft125),
	.ShiftLeft126(ShiftLeft126),
	.ShiftLeft127(ShiftLeft127),
	.ShiftLeft128(ShiftLeft128),
	.ShiftLeft129(ShiftLeft129),
	.ShiftLeft130(ShiftLeft130),
	.ShiftLeft131(ShiftLeft131),
	.ShiftLeft132(ShiftLeft132),
	.ShiftLeft133(ShiftLeft133),
	.ShiftLeft134(ShiftLeft134),
	.ShiftLeft135(ShiftLeft135),
	.ShiftLeft136(ShiftLeft136),
	.ShiftLeft137(ShiftLeft137),
	.ShiftLeft138(ShiftLeft138),
	.ShiftLeft139(ShiftLeft139),
	.ShiftLeft140(ShiftLeft140),
	.ShiftLeft141(ShiftLeft141),
	.ShiftLeft142(ShiftLeft142),
	.ShiftLeft143(ShiftLeft143),
	.ShiftLeft144(ShiftLeft144),
	.ShiftLeft145(ShiftLeft145),
	.ShiftLeft146(ShiftLeft146),
	.ShiftLeft147(ShiftLeft147),
	.ShiftLeft148(ShiftLeft148),
	.ShiftLeft149(ShiftLeft149),
	.ShiftLeft150(ShiftLeft150),
	.ShiftLeft151(ShiftLeft151),
	.ShiftLeft152(ShiftLeft152),
	.ShiftLeft153(ShiftLeft153),
	.ShiftLeft154(ShiftLeft154),
	.ShiftLeft155(ShiftLeft155),
	.ShiftLeft156(ShiftLeft156),
	.ShiftLeft157(ShiftLeft157),
	.ShiftLeft158(ShiftLeft158),
	.ShiftLeft159(ShiftLeft159),
	.ShiftLeft160(ShiftLeft160),
	.ShiftLeft161(ShiftLeft161),
	.ShiftLeft162(ShiftLeft162),
	.ShiftLeft163(ShiftLeft163),
	.ShiftLeft0(ShiftLeft0),
	.ShiftLeft01(ShiftLeft01),
	.ShiftLeft02(ShiftLeft02),
	.ShiftLeft03(ShiftLeft03),
	.ShiftLeft04(ShiftLeft04),
	.ShiftLeft05(ShiftLeft05),
	.ShiftLeft06(ShiftLeft06),
	.ShiftLeft07(ShiftLeft07),
	.reset(altera_reset_synchronizer_int_chain_out),
	.bready(bready1),
	.write_cp_ready(write_cp_ready),
	.src_payload(src_payload1));

cyclonev_lcell_comb arvalid(
	.dataa(!mem_used_7),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(arvalid1),
	.sumout(),
	.cout(),
	.shareout());
defparam arvalid.extended_lut = "off";
defparam arvalid.lut_mask = 64'h2222222222222222;
defparam arvalid.shared_arith = "off";

dffeas address_taken(
	.clk(outclk_wire_0),
	.d(\address_taken~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(address_taken1),
	.prn(vcc));
defparam address_taken.is_wysiwyg = "true";
defparam address_taken.power_up = "low";

cyclonev_lcell_comb awvalid(
	.dataa(!address_taken1),
	.datab(!mem_used_71),
	.datac(!src_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(awvalid1),
	.sumout(),
	.cout(),
	.shareout());
defparam awvalid.extended_lut = "off";
defparam awvalid.lut_mask = 64'h0808080808080808;
defparam awvalid.shared_arith = "off";

cyclonev_lcell_comb \bready~0 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!mem_105_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(bready),
	.sumout(),
	.cout(),
	.shareout());
defparam \bready~0 .extended_lut = "off";
defparam \bready~0 .lut_mask = 64'h1515151515151515;
defparam \bready~0 .shared_arith = "off";

dffeas data_taken(
	.clk(outclk_wire_0),
	.d(\data_taken~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_taken1),
	.prn(vcc));
defparam data_taken.is_wysiwyg = "true";
defparam data_taken.power_up = "low";

cyclonev_lcell_comb wvalid(
	.dataa(!mem_used_71),
	.datab(!src_valid),
	.datac(!data_taken1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wvalid1),
	.sumout(),
	.cout(),
	.shareout());
defparam wvalid.extended_lut = "off";
defparam wvalid.lut_mask = 64'h2020202020202020;
defparam wvalid.shared_arith = "off";

cyclonev_lcell_comb \bready~1 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(bready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \bready~1 .extended_lut = "off";
defparam \bready~1 .lut_mask = 64'h1111111111111111;
defparam \bready~1 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_ready~0 (
	.dataa(!f2h_AWREADY_0),
	.datab(!f2h_WREADY_0),
	.datac(!address_taken1),
	.datad(!mem_used_71),
	.datae(!data_taken1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_ready~0 .extended_lut = "off";
defparam \write_cp_ready~0 .lut_mask = 64'h1303575713035757;
defparam \write_cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \address_taken~0 (
	.dataa(!f2h_AWREADY_0),
	.datab(!address_taken1),
	.datac(!awvalid1),
	.datad(!fifo_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_taken~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_taken~0 .extended_lut = "off";
defparam \address_taken~0 .lut_mask = 64'h3700370037003700;
defparam \address_taken~0 .shared_arith = "off";

cyclonev_lcell_comb \data_taken~0 (
	.dataa(!f2h_WREADY_0),
	.datab(!data_taken1),
	.datac(!wvalid1),
	.datad(!fifo_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_taken~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_taken~0 .extended_lut = "off";
defparam \data_taken~0 .lut_mask = 64'h3700370037003700;
defparam \data_taken~0 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_4 (
	f2h_ARREADY_0,
	f2h_RVALID_0,
	clk,
	mem_113_0,
	mem_68_0,
	mem_64_0,
	mem_used_7,
	saved_grant_0,
	last_channel_1,
	has_pending_responses,
	read_select,
	hold_waitrequest,
	write,
	src_payload,
	reset,
	ShiftLeft0)/* synthesis synthesis_greybox=0 */;
input 	f2h_ARREADY_0;
input 	f2h_RVALID_0;
input 	clk;
output 	mem_113_0;
output 	mem_68_0;
output 	mem_64_0;
output 	mem_used_7;
input 	saved_grant_0;
input 	last_channel_1;
input 	has_pending_responses;
input 	read_select;
input 	hold_waitrequest;
output 	write;
input 	src_payload;
input 	reset;
input 	ShiftLeft0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[7][154]~q ;
wire \mem~0_combout ;
wire \write~1_combout ;
wire \mem_used~2_combout ;
wire \mem_used[6]~3_combout ;
wire \mem_used[6]~q ;
wire \mem_used~5_combout ;
wire \mem_used[5]~q ;
wire \mem_used~7_combout ;
wire \mem_used[4]~q ;
wire \mem_used~8_combout ;
wire \mem_used[3]~q ;
wire \mem_used~6_combout ;
wire \mem_used[2]~q ;
wire \mem_used~4_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \always6~0_combout ;
wire \mem[6][113]~q ;
wire \always5~0_combout ;
wire \mem[5][113]~q ;
wire \always4~0_combout ;
wire \mem[4][113]~q ;
wire \always3~0_combout ;
wire \mem[3][113]~q ;
wire \always2~0_combout ;
wire \mem[2][113]~q ;
wire \always1~0_combout ;
wire \mem[1][113]~q ;
wire \always0~0_combout ;
wire \mem[7][68]~q ;
wire \mem~1_combout ;
wire \mem[6][68]~q ;
wire \mem[5][68]~q ;
wire \mem[4][68]~q ;
wire \mem[3][68]~q ;
wire \mem[2][68]~q ;
wire \mem[1][68]~q ;
wire \mem[7][64]~q ;
wire \mem~2_combout ;
wire \mem[6][64]~q ;
wire \mem[5][64]~q ;
wire \mem[4][64]~q ;
wire \mem[3][64]~q ;
wire \mem[2][64]~q ;
wire \mem[1][64]~q ;
wire \mem_used[7]~0_combout ;


dffeas \mem[0][113] (
	.clk(clk),
	.d(saved_grant_0),
	.asdata(\mem[1][113]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[1][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[1][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_64_0),
	.prn(vcc));
defparam \mem[0][64] .is_wysiwyg = "true";
defparam \mem[0][64] .power_up = "low";

dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used[7]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_7),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!saved_grant_0),
	.datab(!last_channel_1),
	.datac(!has_pending_responses),
	.datad(!read_select),
	.datae(!hold_waitrequest),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0000005100000051;
defparam \write~0 .shared_arith = "off";

dffeas \mem[7][154] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][154]~q ),
	.prn(vcc));
defparam \mem[7][154] .is_wysiwyg = "true";
defparam \mem[7][154] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_7),
	.datab(!saved_grant_0),
	.datac(!\mem[7][154]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!f2h_ARREADY_0),
	.datab(!mem_used_7),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0404040404040404;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used~2 (
	.dataa(!mem_used_7),
	.datab(!\write~1_combout ),
	.datac(!\mem_used[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~2 .extended_lut = "off";
defparam \mem_used~2 .lut_mask = 64'h5757575757575757;
defparam \mem_used~2 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[6]~3 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\write~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[6]~3 .extended_lut = "off";
defparam \mem_used[6]~3 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \mem_used[6]~3 .shared_arith = "off";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cyclonev_lcell_comb \mem_used~5 (
	.dataa(!\write~1_combout ),
	.datab(!\mem_used[6]~q ),
	.datac(!\mem_used[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~5 .extended_lut = "off";
defparam \mem_used~5 .lut_mask = 64'h2727272727272727;
defparam \mem_used~5 .shared_arith = "off";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cyclonev_lcell_comb \mem_used~7 (
	.dataa(!\write~1_combout ),
	.datab(!\mem_used[5]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~7 .extended_lut = "off";
defparam \mem_used~7 .lut_mask = 64'h2727272727272727;
defparam \mem_used~7 .shared_arith = "off";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cyclonev_lcell_comb \mem_used~8 (
	.dataa(!\write~1_combout ),
	.datab(!\mem_used[2]~q ),
	.datac(!\mem_used[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~8 .extended_lut = "off";
defparam \mem_used~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_used~8 .shared_arith = "off";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cyclonev_lcell_comb \mem_used~6 (
	.dataa(!\write~1_combout ),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~6 .extended_lut = "off";
defparam \mem_used~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_used~6 .shared_arith = "off";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cyclonev_lcell_comb \mem_used~4 (
	.dataa(!\mem_used[0]~q ),
	.datab(!\write~1_combout ),
	.datac(!\mem_used[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~4 .extended_lut = "off";
defparam \mem_used~4 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \mem_used~4 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\write~1_combout ),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h2F3F2F3F2F3F2F3F;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always6~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \always6~0 .shared_arith = "off";

dffeas \mem[6][113] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][113]~q ),
	.prn(vcc));
defparam \mem[6][113] .is_wysiwyg = "true";
defparam \mem[6][113] .power_up = "low";

cyclonev_lcell_comb \always5~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \always5~0 .shared_arith = "off";

dffeas \mem[5][113] (
	.clk(clk),
	.d(saved_grant_0),
	.asdata(\mem[6][113]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][113]~q ),
	.prn(vcc));
defparam \mem[5][113] .is_wysiwyg = "true";
defparam \mem[5][113] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[4][113] (
	.clk(clk),
	.d(saved_grant_0),
	.asdata(\mem[5][113]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][113]~q ),
	.prn(vcc));
defparam \mem[4][113] .is_wysiwyg = "true";
defparam \mem[4][113] .power_up = "low";

cyclonev_lcell_comb \always3~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \always3~0 .shared_arith = "off";

dffeas \mem[3][113] (
	.clk(clk),
	.d(saved_grant_0),
	.asdata(\mem[4][113]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][113]~q ),
	.prn(vcc));
defparam \mem[3][113] .is_wysiwyg = "true";
defparam \mem[3][113] .power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \always2~0 .shared_arith = "off";

dffeas \mem[2][113] (
	.clk(clk),
	.d(saved_grant_0),
	.asdata(\mem[3][113]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][113]~q ),
	.prn(vcc));
defparam \mem[2][113] .is_wysiwyg = "true";
defparam \mem[2][113] .power_up = "low";

cyclonev_lcell_comb \always1~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(!\mem_used[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \always1~0 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(saved_grant_0),
	.asdata(\mem[2][113]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[7][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][68]~q ),
	.prn(vcc));
defparam \mem[7][68] .is_wysiwyg = "true";
defparam \mem[7][68] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_7),
	.datab(!src_payload),
	.datac(!\mem[7][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[6][68] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][68]~q ),
	.prn(vcc));
defparam \mem[6][68] .is_wysiwyg = "true";
defparam \mem[6][68] .power_up = "low";

dffeas \mem[5][68] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[6][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][68]~q ),
	.prn(vcc));
defparam \mem[5][68] .is_wysiwyg = "true";
defparam \mem[5][68] .power_up = "low";

dffeas \mem[4][68] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[5][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][68]~q ),
	.prn(vcc));
defparam \mem[4][68] .is_wysiwyg = "true";
defparam \mem[4][68] .power_up = "low";

dffeas \mem[3][68] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[4][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][68]~q ),
	.prn(vcc));
defparam \mem[3][68] .is_wysiwyg = "true";
defparam \mem[3][68] .power_up = "low";

dffeas \mem[2][68] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[3][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][68]~q ),
	.prn(vcc));
defparam \mem[2][68] .is_wysiwyg = "true";
defparam \mem[2][68] .power_up = "low";

dffeas \mem[1][68] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[2][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

dffeas \mem[7][64] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][64]~q ),
	.prn(vcc));
defparam \mem[7][64] .is_wysiwyg = "true";
defparam \mem[7][64] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft0),
	.datac(!\mem[7][64]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[6][64] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][64]~q ),
	.prn(vcc));
defparam \mem[6][64] .is_wysiwyg = "true";
defparam \mem[6][64] .power_up = "low";

dffeas \mem[5][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[6][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][64]~q ),
	.prn(vcc));
defparam \mem[5][64] .is_wysiwyg = "true";
defparam \mem[5][64] .power_up = "low";

dffeas \mem[4][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[5][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][64]~q ),
	.prn(vcc));
defparam \mem[4][64] .is_wysiwyg = "true";
defparam \mem[4][64] .power_up = "low";

dffeas \mem[3][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[4][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][64]~q ),
	.prn(vcc));
defparam \mem[3][64] .is_wysiwyg = "true";
defparam \mem[3][64] .power_up = "low";

dffeas \mem[2][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[3][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][64]~q ),
	.prn(vcc));
defparam \mem[2][64] .is_wysiwyg = "true";
defparam \mem[2][64] .power_up = "low";

dffeas \mem[1][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[2][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][64]~q ),
	.prn(vcc));
defparam \mem[1][64] .is_wysiwyg = "true";
defparam \mem[1][64] .power_up = "low";

cyclonev_lcell_comb \mem_used[7]~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!mem_used_7),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~1_combout ),
	.datae(!\mem_used[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[7]~0 .extended_lut = "off";
defparam \mem_used[7]~0 .lut_mask = 64'h320132FB320132FB;
defparam \mem_used[7]~0 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_5 (
	f2h_BVALID_0,
	clk,
	mem_105_0,
	mem_139_0,
	mem_68_0,
	mem_64_0,
	mem_69_0,
	mem_65_0,
	mem_70_0,
	mem_66_0,
	mem_71_0,
	mem_67_0,
	mem_8_0,
	mem_40_0,
	mem_16_0,
	mem_48_0,
	mem_24_0,
	mem_56_0,
	mem_0_0,
	mem_32_0,
	mem_9_0,
	mem_41_0,
	mem_17_0,
	mem_49_0,
	mem_25_0,
	mem_57_0,
	mem_1_0,
	mem_33_0,
	mem_10_0,
	mem_42_0,
	mem_18_0,
	mem_50_0,
	mem_26_0,
	mem_58_0,
	mem_2_0,
	mem_34_0,
	mem_11_0,
	mem_43_0,
	mem_19_0,
	mem_51_0,
	mem_27_0,
	mem_59_0,
	mem_3_0,
	mem_35_0,
	mem_12_0,
	mem_44_0,
	mem_20_0,
	mem_52_0,
	mem_28_0,
	mem_60_0,
	mem_4_0,
	mem_36_0,
	mem_13_0,
	mem_45_0,
	mem_21_0,
	mem_53_0,
	mem_29_0,
	mem_61_0,
	mem_5_0,
	mem_37_0,
	mem_14_0,
	mem_46_0,
	mem_22_0,
	mem_54_0,
	mem_30_0,
	mem_62_0,
	mem_6_0,
	mem_38_0,
	mem_15_0,
	mem_47_0,
	mem_23_0,
	mem_55_0,
	mem_31_0,
	mem_63_0,
	mem_7_0,
	mem_39_0,
	mem_used_7,
	saved_grant_1,
	src_valid,
	mem_used_0,
	ShiftLeft1,
	ShiftLeft11,
	ShiftLeft12,
	ShiftLeft13,
	ShiftLeft14,
	ShiftLeft15,
	ShiftLeft16,
	ShiftLeft17,
	ShiftLeft18,
	ShiftLeft19,
	ShiftLeft110,
	ShiftLeft111,
	ShiftLeft112,
	ShiftLeft113,
	ShiftLeft114,
	ShiftLeft115,
	ShiftLeft116,
	ShiftLeft117,
	ShiftLeft118,
	ShiftLeft119,
	ShiftLeft120,
	ShiftLeft121,
	ShiftLeft122,
	ShiftLeft123,
	ShiftLeft124,
	ShiftLeft125,
	ShiftLeft126,
	ShiftLeft127,
	ShiftLeft128,
	ShiftLeft129,
	ShiftLeft130,
	ShiftLeft131,
	ShiftLeft132,
	ShiftLeft133,
	ShiftLeft134,
	ShiftLeft135,
	ShiftLeft136,
	ShiftLeft137,
	ShiftLeft138,
	ShiftLeft139,
	ShiftLeft140,
	ShiftLeft141,
	ShiftLeft142,
	ShiftLeft143,
	ShiftLeft144,
	ShiftLeft145,
	ShiftLeft146,
	ShiftLeft147,
	ShiftLeft148,
	ShiftLeft149,
	ShiftLeft150,
	ShiftLeft151,
	ShiftLeft152,
	ShiftLeft153,
	ShiftLeft154,
	ShiftLeft155,
	ShiftLeft156,
	ShiftLeft157,
	ShiftLeft158,
	ShiftLeft159,
	ShiftLeft160,
	ShiftLeft161,
	ShiftLeft162,
	ShiftLeft163,
	ShiftLeft0,
	ShiftLeft01,
	ShiftLeft02,
	ShiftLeft03,
	ShiftLeft04,
	ShiftLeft05,
	ShiftLeft06,
	ShiftLeft07,
	reset,
	bready,
	write_cp_ready,
	src_payload)/* synthesis synthesis_greybox=0 */;
input 	f2h_BVALID_0;
input 	clk;
output 	mem_105_0;
output 	mem_139_0;
output 	mem_68_0;
output 	mem_64_0;
output 	mem_69_0;
output 	mem_65_0;
output 	mem_70_0;
output 	mem_66_0;
output 	mem_71_0;
output 	mem_67_0;
output 	mem_8_0;
output 	mem_40_0;
output 	mem_16_0;
output 	mem_48_0;
output 	mem_24_0;
output 	mem_56_0;
output 	mem_0_0;
output 	mem_32_0;
output 	mem_9_0;
output 	mem_41_0;
output 	mem_17_0;
output 	mem_49_0;
output 	mem_25_0;
output 	mem_57_0;
output 	mem_1_0;
output 	mem_33_0;
output 	mem_10_0;
output 	mem_42_0;
output 	mem_18_0;
output 	mem_50_0;
output 	mem_26_0;
output 	mem_58_0;
output 	mem_2_0;
output 	mem_34_0;
output 	mem_11_0;
output 	mem_43_0;
output 	mem_19_0;
output 	mem_51_0;
output 	mem_27_0;
output 	mem_59_0;
output 	mem_3_0;
output 	mem_35_0;
output 	mem_12_0;
output 	mem_44_0;
output 	mem_20_0;
output 	mem_52_0;
output 	mem_28_0;
output 	mem_60_0;
output 	mem_4_0;
output 	mem_36_0;
output 	mem_13_0;
output 	mem_45_0;
output 	mem_21_0;
output 	mem_53_0;
output 	mem_29_0;
output 	mem_61_0;
output 	mem_5_0;
output 	mem_37_0;
output 	mem_14_0;
output 	mem_46_0;
output 	mem_22_0;
output 	mem_54_0;
output 	mem_30_0;
output 	mem_62_0;
output 	mem_6_0;
output 	mem_38_0;
output 	mem_15_0;
output 	mem_47_0;
output 	mem_23_0;
output 	mem_55_0;
output 	mem_31_0;
output 	mem_63_0;
output 	mem_7_0;
output 	mem_39_0;
output 	mem_used_7;
input 	saved_grant_1;
input 	src_valid;
output 	mem_used_0;
input 	ShiftLeft1;
input 	ShiftLeft11;
input 	ShiftLeft12;
input 	ShiftLeft13;
input 	ShiftLeft14;
input 	ShiftLeft15;
input 	ShiftLeft16;
input 	ShiftLeft17;
input 	ShiftLeft18;
input 	ShiftLeft19;
input 	ShiftLeft110;
input 	ShiftLeft111;
input 	ShiftLeft112;
input 	ShiftLeft113;
input 	ShiftLeft114;
input 	ShiftLeft115;
input 	ShiftLeft116;
input 	ShiftLeft117;
input 	ShiftLeft118;
input 	ShiftLeft119;
input 	ShiftLeft120;
input 	ShiftLeft121;
input 	ShiftLeft122;
input 	ShiftLeft123;
input 	ShiftLeft124;
input 	ShiftLeft125;
input 	ShiftLeft126;
input 	ShiftLeft127;
input 	ShiftLeft128;
input 	ShiftLeft129;
input 	ShiftLeft130;
input 	ShiftLeft131;
input 	ShiftLeft132;
input 	ShiftLeft133;
input 	ShiftLeft134;
input 	ShiftLeft135;
input 	ShiftLeft136;
input 	ShiftLeft137;
input 	ShiftLeft138;
input 	ShiftLeft139;
input 	ShiftLeft140;
input 	ShiftLeft141;
input 	ShiftLeft142;
input 	ShiftLeft143;
input 	ShiftLeft144;
input 	ShiftLeft145;
input 	ShiftLeft146;
input 	ShiftLeft147;
input 	ShiftLeft148;
input 	ShiftLeft149;
input 	ShiftLeft150;
input 	ShiftLeft151;
input 	ShiftLeft152;
input 	ShiftLeft153;
input 	ShiftLeft154;
input 	ShiftLeft155;
input 	ShiftLeft156;
input 	ShiftLeft157;
input 	ShiftLeft158;
input 	ShiftLeft159;
input 	ShiftLeft160;
input 	ShiftLeft161;
input 	ShiftLeft162;
input 	ShiftLeft163;
input 	ShiftLeft0;
input 	ShiftLeft01;
input 	ShiftLeft02;
input 	ShiftLeft03;
input 	ShiftLeft04;
input 	ShiftLeft05;
input 	ShiftLeft06;
input 	ShiftLeft07;
input 	reset;
input 	bready;
input 	write_cp_ready;
input 	src_payload;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[7][106]~q ;
wire \mem~0_combout ;
wire \write~0_combout ;
wire \mem_used~4_combout ;
wire \mem_used[6]~3_combout ;
wire \mem_used[1]~q ;
wire \mem_used~6_combout ;
wire \mem_used[2]~q ;
wire \mem_used~8_combout ;
wire \mem_used[3]~q ;
wire \mem_used~7_combout ;
wire \mem_used[4]~q ;
wire \mem_used~5_combout ;
wire \mem_used[5]~q ;
wire \mem_used~2_combout ;
wire \mem_used[6]~q ;
wire \always6~0_combout ;
wire \mem[6][105]~q ;
wire \always5~0_combout ;
wire \mem[5][105]~q ;
wire \always4~0_combout ;
wire \mem[4][105]~q ;
wire \always3~0_combout ;
wire \mem[3][105]~q ;
wire \always2~0_combout ;
wire \mem[2][105]~q ;
wire \always1~0_combout ;
wire \mem[1][105]~q ;
wire \always0~0_combout ;
wire \mem[7][154]~q ;
wire \mem~1_combout ;
wire \mem[6][139]~q ;
wire \mem[5][139]~q ;
wire \mem[4][139]~q ;
wire \mem[3][139]~q ;
wire \mem[2][139]~q ;
wire \mem[1][139]~q ;
wire \mem[7][68]~q ;
wire \mem~2_combout ;
wire \mem[6][68]~q ;
wire \mem[5][68]~q ;
wire \mem[4][68]~q ;
wire \mem[3][68]~q ;
wire \mem[2][68]~q ;
wire \mem[1][68]~q ;
wire \mem[7][64]~q ;
wire \mem~3_combout ;
wire \mem[6][64]~q ;
wire \mem[5][64]~q ;
wire \mem[4][64]~q ;
wire \mem[3][64]~q ;
wire \mem[2][64]~q ;
wire \mem[1][64]~q ;
wire \mem[7][69]~q ;
wire \mem~4_combout ;
wire \mem[6][69]~q ;
wire \mem[5][69]~q ;
wire \mem[4][69]~q ;
wire \mem[3][69]~q ;
wire \mem[2][69]~q ;
wire \mem[1][69]~q ;
wire \mem[7][65]~q ;
wire \mem~5_combout ;
wire \mem[6][65]~q ;
wire \mem[5][65]~q ;
wire \mem[4][65]~q ;
wire \mem[3][65]~q ;
wire \mem[2][65]~q ;
wire \mem[1][65]~q ;
wire \mem[7][70]~q ;
wire \mem~6_combout ;
wire \mem[6][70]~q ;
wire \mem[5][70]~q ;
wire \mem[4][70]~q ;
wire \mem[3][70]~q ;
wire \mem[2][70]~q ;
wire \mem[1][70]~q ;
wire \mem[7][66]~q ;
wire \mem~7_combout ;
wire \mem[6][66]~q ;
wire \mem[5][66]~q ;
wire \mem[4][66]~q ;
wire \mem[3][66]~q ;
wire \mem[2][66]~q ;
wire \mem[1][66]~q ;
wire \mem[7][71]~q ;
wire \mem~8_combout ;
wire \mem[6][71]~q ;
wire \mem[5][71]~q ;
wire \mem[4][71]~q ;
wire \mem[3][71]~q ;
wire \mem[2][71]~q ;
wire \mem[1][71]~q ;
wire \mem[7][67]~q ;
wire \mem~9_combout ;
wire \mem[6][67]~q ;
wire \mem[5][67]~q ;
wire \mem[4][67]~q ;
wire \mem[3][67]~q ;
wire \mem[2][67]~q ;
wire \mem[1][67]~q ;
wire \mem[7][8]~q ;
wire \mem~10_combout ;
wire \mem[6][8]~q ;
wire \mem[5][8]~q ;
wire \mem[4][8]~q ;
wire \mem[3][8]~q ;
wire \mem[2][8]~q ;
wire \mem[1][8]~q ;
wire \mem[7][40]~q ;
wire \mem~11_combout ;
wire \mem[6][40]~q ;
wire \mem[5][40]~q ;
wire \mem[4][40]~q ;
wire \mem[3][40]~q ;
wire \mem[2][40]~q ;
wire \mem[1][40]~q ;
wire \mem[7][16]~q ;
wire \mem~12_combout ;
wire \mem[6][16]~q ;
wire \mem[5][16]~q ;
wire \mem[4][16]~q ;
wire \mem[3][16]~q ;
wire \mem[2][16]~q ;
wire \mem[1][16]~q ;
wire \mem[7][48]~q ;
wire \mem~13_combout ;
wire \mem[6][48]~q ;
wire \mem[5][48]~q ;
wire \mem[4][48]~q ;
wire \mem[3][48]~q ;
wire \mem[2][48]~q ;
wire \mem[1][48]~q ;
wire \mem[7][24]~q ;
wire \mem~14_combout ;
wire \mem[6][24]~q ;
wire \mem[5][24]~q ;
wire \mem[4][24]~q ;
wire \mem[3][24]~q ;
wire \mem[2][24]~q ;
wire \mem[1][24]~q ;
wire \mem[7][56]~q ;
wire \mem~15_combout ;
wire \mem[6][56]~q ;
wire \mem[5][56]~q ;
wire \mem[4][56]~q ;
wire \mem[3][56]~q ;
wire \mem[2][56]~q ;
wire \mem[1][56]~q ;
wire \mem[7][0]~q ;
wire \mem~16_combout ;
wire \mem[6][0]~q ;
wire \mem[5][0]~q ;
wire \mem[4][0]~q ;
wire \mem[3][0]~q ;
wire \mem[2][0]~q ;
wire \mem[1][0]~q ;
wire \mem[7][32]~q ;
wire \mem~17_combout ;
wire \mem[6][32]~q ;
wire \mem[5][32]~q ;
wire \mem[4][32]~q ;
wire \mem[3][32]~q ;
wire \mem[2][32]~q ;
wire \mem[1][32]~q ;
wire \mem[7][9]~q ;
wire \mem~18_combout ;
wire \mem[6][9]~q ;
wire \mem[5][9]~q ;
wire \mem[4][9]~q ;
wire \mem[3][9]~q ;
wire \mem[2][9]~q ;
wire \mem[1][9]~q ;
wire \mem[7][41]~q ;
wire \mem~19_combout ;
wire \mem[6][41]~q ;
wire \mem[5][41]~q ;
wire \mem[4][41]~q ;
wire \mem[3][41]~q ;
wire \mem[2][41]~q ;
wire \mem[1][41]~q ;
wire \mem[7][17]~q ;
wire \mem~20_combout ;
wire \mem[6][17]~q ;
wire \mem[5][17]~q ;
wire \mem[4][17]~q ;
wire \mem[3][17]~q ;
wire \mem[2][17]~q ;
wire \mem[1][17]~q ;
wire \mem[7][49]~q ;
wire \mem~21_combout ;
wire \mem[6][49]~q ;
wire \mem[5][49]~q ;
wire \mem[4][49]~q ;
wire \mem[3][49]~q ;
wire \mem[2][49]~q ;
wire \mem[1][49]~q ;
wire \mem[7][25]~q ;
wire \mem~22_combout ;
wire \mem[6][25]~q ;
wire \mem[5][25]~q ;
wire \mem[4][25]~q ;
wire \mem[3][25]~q ;
wire \mem[2][25]~q ;
wire \mem[1][25]~q ;
wire \mem[7][57]~q ;
wire \mem~23_combout ;
wire \mem[6][57]~q ;
wire \mem[5][57]~q ;
wire \mem[4][57]~q ;
wire \mem[3][57]~q ;
wire \mem[2][57]~q ;
wire \mem[1][57]~q ;
wire \mem[7][1]~q ;
wire \mem~24_combout ;
wire \mem[6][1]~q ;
wire \mem[5][1]~q ;
wire \mem[4][1]~q ;
wire \mem[3][1]~q ;
wire \mem[2][1]~q ;
wire \mem[1][1]~q ;
wire \mem[7][33]~q ;
wire \mem~25_combout ;
wire \mem[6][33]~q ;
wire \mem[5][33]~q ;
wire \mem[4][33]~q ;
wire \mem[3][33]~q ;
wire \mem[2][33]~q ;
wire \mem[1][33]~q ;
wire \mem[7][10]~q ;
wire \mem~26_combout ;
wire \mem[6][10]~q ;
wire \mem[5][10]~q ;
wire \mem[4][10]~q ;
wire \mem[3][10]~q ;
wire \mem[2][10]~q ;
wire \mem[1][10]~q ;
wire \mem[7][42]~q ;
wire \mem~27_combout ;
wire \mem[6][42]~q ;
wire \mem[5][42]~q ;
wire \mem[4][42]~q ;
wire \mem[3][42]~q ;
wire \mem[2][42]~q ;
wire \mem[1][42]~q ;
wire \mem[7][18]~q ;
wire \mem~28_combout ;
wire \mem[6][18]~q ;
wire \mem[5][18]~q ;
wire \mem[4][18]~q ;
wire \mem[3][18]~q ;
wire \mem[2][18]~q ;
wire \mem[1][18]~q ;
wire \mem[7][50]~q ;
wire \mem~29_combout ;
wire \mem[6][50]~q ;
wire \mem[5][50]~q ;
wire \mem[4][50]~q ;
wire \mem[3][50]~q ;
wire \mem[2][50]~q ;
wire \mem[1][50]~q ;
wire \mem[7][26]~q ;
wire \mem~30_combout ;
wire \mem[6][26]~q ;
wire \mem[5][26]~q ;
wire \mem[4][26]~q ;
wire \mem[3][26]~q ;
wire \mem[2][26]~q ;
wire \mem[1][26]~q ;
wire \mem[7][58]~q ;
wire \mem~31_combout ;
wire \mem[6][58]~q ;
wire \mem[5][58]~q ;
wire \mem[4][58]~q ;
wire \mem[3][58]~q ;
wire \mem[2][58]~q ;
wire \mem[1][58]~q ;
wire \mem[7][2]~q ;
wire \mem~32_combout ;
wire \mem[6][2]~q ;
wire \mem[5][2]~q ;
wire \mem[4][2]~q ;
wire \mem[3][2]~q ;
wire \mem[2][2]~q ;
wire \mem[1][2]~q ;
wire \mem[7][34]~q ;
wire \mem~33_combout ;
wire \mem[6][34]~q ;
wire \mem[5][34]~q ;
wire \mem[4][34]~q ;
wire \mem[3][34]~q ;
wire \mem[2][34]~q ;
wire \mem[1][34]~q ;
wire \mem[7][11]~q ;
wire \mem~34_combout ;
wire \mem[6][11]~q ;
wire \mem[5][11]~q ;
wire \mem[4][11]~q ;
wire \mem[3][11]~q ;
wire \mem[2][11]~q ;
wire \mem[1][11]~q ;
wire \mem[7][43]~q ;
wire \mem~35_combout ;
wire \mem[6][43]~q ;
wire \mem[5][43]~q ;
wire \mem[4][43]~q ;
wire \mem[3][43]~q ;
wire \mem[2][43]~q ;
wire \mem[1][43]~q ;
wire \mem[7][19]~q ;
wire \mem~36_combout ;
wire \mem[6][19]~q ;
wire \mem[5][19]~q ;
wire \mem[4][19]~q ;
wire \mem[3][19]~q ;
wire \mem[2][19]~q ;
wire \mem[1][19]~q ;
wire \mem[7][51]~q ;
wire \mem~37_combout ;
wire \mem[6][51]~q ;
wire \mem[5][51]~q ;
wire \mem[4][51]~q ;
wire \mem[3][51]~q ;
wire \mem[2][51]~q ;
wire \mem[1][51]~q ;
wire \mem[7][27]~q ;
wire \mem~38_combout ;
wire \mem[6][27]~q ;
wire \mem[5][27]~q ;
wire \mem[4][27]~q ;
wire \mem[3][27]~q ;
wire \mem[2][27]~q ;
wire \mem[1][27]~q ;
wire \mem[7][59]~q ;
wire \mem~39_combout ;
wire \mem[6][59]~q ;
wire \mem[5][59]~q ;
wire \mem[4][59]~q ;
wire \mem[3][59]~q ;
wire \mem[2][59]~q ;
wire \mem[1][59]~q ;
wire \mem[7][3]~q ;
wire \mem~40_combout ;
wire \mem[6][3]~q ;
wire \mem[5][3]~q ;
wire \mem[4][3]~q ;
wire \mem[3][3]~q ;
wire \mem[2][3]~q ;
wire \mem[1][3]~q ;
wire \mem[7][35]~q ;
wire \mem~41_combout ;
wire \mem[6][35]~q ;
wire \mem[5][35]~q ;
wire \mem[4][35]~q ;
wire \mem[3][35]~q ;
wire \mem[2][35]~q ;
wire \mem[1][35]~q ;
wire \mem[7][12]~q ;
wire \mem~42_combout ;
wire \mem[6][12]~q ;
wire \mem[5][12]~q ;
wire \mem[4][12]~q ;
wire \mem[3][12]~q ;
wire \mem[2][12]~q ;
wire \mem[1][12]~q ;
wire \mem[7][44]~q ;
wire \mem~43_combout ;
wire \mem[6][44]~q ;
wire \mem[5][44]~q ;
wire \mem[4][44]~q ;
wire \mem[3][44]~q ;
wire \mem[2][44]~q ;
wire \mem[1][44]~q ;
wire \mem[7][20]~q ;
wire \mem~44_combout ;
wire \mem[6][20]~q ;
wire \mem[5][20]~q ;
wire \mem[4][20]~q ;
wire \mem[3][20]~q ;
wire \mem[2][20]~q ;
wire \mem[1][20]~q ;
wire \mem[7][52]~q ;
wire \mem~45_combout ;
wire \mem[6][52]~q ;
wire \mem[5][52]~q ;
wire \mem[4][52]~q ;
wire \mem[3][52]~q ;
wire \mem[2][52]~q ;
wire \mem[1][52]~q ;
wire \mem[7][28]~q ;
wire \mem~46_combout ;
wire \mem[6][28]~q ;
wire \mem[5][28]~q ;
wire \mem[4][28]~q ;
wire \mem[3][28]~q ;
wire \mem[2][28]~q ;
wire \mem[1][28]~q ;
wire \mem[7][60]~q ;
wire \mem~47_combout ;
wire \mem[6][60]~q ;
wire \mem[5][60]~q ;
wire \mem[4][60]~q ;
wire \mem[3][60]~q ;
wire \mem[2][60]~q ;
wire \mem[1][60]~q ;
wire \mem[7][4]~q ;
wire \mem~48_combout ;
wire \mem[6][4]~q ;
wire \mem[5][4]~q ;
wire \mem[4][4]~q ;
wire \mem[3][4]~q ;
wire \mem[2][4]~q ;
wire \mem[1][4]~q ;
wire \mem[7][36]~q ;
wire \mem~49_combout ;
wire \mem[6][36]~q ;
wire \mem[5][36]~q ;
wire \mem[4][36]~q ;
wire \mem[3][36]~q ;
wire \mem[2][36]~q ;
wire \mem[1][36]~q ;
wire \mem[7][13]~q ;
wire \mem~50_combout ;
wire \mem[6][13]~q ;
wire \mem[5][13]~q ;
wire \mem[4][13]~q ;
wire \mem[3][13]~q ;
wire \mem[2][13]~q ;
wire \mem[1][13]~q ;
wire \mem[7][45]~q ;
wire \mem~51_combout ;
wire \mem[6][45]~q ;
wire \mem[5][45]~q ;
wire \mem[4][45]~q ;
wire \mem[3][45]~q ;
wire \mem[2][45]~q ;
wire \mem[1][45]~q ;
wire \mem[7][21]~q ;
wire \mem~52_combout ;
wire \mem[6][21]~q ;
wire \mem[5][21]~q ;
wire \mem[4][21]~q ;
wire \mem[3][21]~q ;
wire \mem[2][21]~q ;
wire \mem[1][21]~q ;
wire \mem[7][53]~q ;
wire \mem~53_combout ;
wire \mem[6][53]~q ;
wire \mem[5][53]~q ;
wire \mem[4][53]~q ;
wire \mem[3][53]~q ;
wire \mem[2][53]~q ;
wire \mem[1][53]~q ;
wire \mem[7][29]~q ;
wire \mem~54_combout ;
wire \mem[6][29]~q ;
wire \mem[5][29]~q ;
wire \mem[4][29]~q ;
wire \mem[3][29]~q ;
wire \mem[2][29]~q ;
wire \mem[1][29]~q ;
wire \mem[7][61]~q ;
wire \mem~55_combout ;
wire \mem[6][61]~q ;
wire \mem[5][61]~q ;
wire \mem[4][61]~q ;
wire \mem[3][61]~q ;
wire \mem[2][61]~q ;
wire \mem[1][61]~q ;
wire \mem[7][5]~q ;
wire \mem~56_combout ;
wire \mem[6][5]~q ;
wire \mem[5][5]~q ;
wire \mem[4][5]~q ;
wire \mem[3][5]~q ;
wire \mem[2][5]~q ;
wire \mem[1][5]~q ;
wire \mem[7][37]~q ;
wire \mem~57_combout ;
wire \mem[6][37]~q ;
wire \mem[5][37]~q ;
wire \mem[4][37]~q ;
wire \mem[3][37]~q ;
wire \mem[2][37]~q ;
wire \mem[1][37]~q ;
wire \mem[7][14]~q ;
wire \mem~58_combout ;
wire \mem[6][14]~q ;
wire \mem[5][14]~q ;
wire \mem[4][14]~q ;
wire \mem[3][14]~q ;
wire \mem[2][14]~q ;
wire \mem[1][14]~q ;
wire \mem[7][46]~q ;
wire \mem~59_combout ;
wire \mem[6][46]~q ;
wire \mem[5][46]~q ;
wire \mem[4][46]~q ;
wire \mem[3][46]~q ;
wire \mem[2][46]~q ;
wire \mem[1][46]~q ;
wire \mem[7][22]~q ;
wire \mem~60_combout ;
wire \mem[6][22]~q ;
wire \mem[5][22]~q ;
wire \mem[4][22]~q ;
wire \mem[3][22]~q ;
wire \mem[2][22]~q ;
wire \mem[1][22]~q ;
wire \mem[7][54]~q ;
wire \mem~61_combout ;
wire \mem[6][54]~q ;
wire \mem[5][54]~q ;
wire \mem[4][54]~q ;
wire \mem[3][54]~q ;
wire \mem[2][54]~q ;
wire \mem[1][54]~q ;
wire \mem[7][30]~q ;
wire \mem~62_combout ;
wire \mem[6][30]~q ;
wire \mem[5][30]~q ;
wire \mem[4][30]~q ;
wire \mem[3][30]~q ;
wire \mem[2][30]~q ;
wire \mem[1][30]~q ;
wire \mem[7][62]~q ;
wire \mem~63_combout ;
wire \mem[6][62]~q ;
wire \mem[5][62]~q ;
wire \mem[4][62]~q ;
wire \mem[3][62]~q ;
wire \mem[2][62]~q ;
wire \mem[1][62]~q ;
wire \mem[7][6]~q ;
wire \mem~64_combout ;
wire \mem[6][6]~q ;
wire \mem[5][6]~q ;
wire \mem[4][6]~q ;
wire \mem[3][6]~q ;
wire \mem[2][6]~q ;
wire \mem[1][6]~q ;
wire \mem[7][38]~q ;
wire \mem~65_combout ;
wire \mem[6][38]~q ;
wire \mem[5][38]~q ;
wire \mem[4][38]~q ;
wire \mem[3][38]~q ;
wire \mem[2][38]~q ;
wire \mem[1][38]~q ;
wire \mem[7][15]~q ;
wire \mem~66_combout ;
wire \mem[6][15]~q ;
wire \mem[5][15]~q ;
wire \mem[4][15]~q ;
wire \mem[3][15]~q ;
wire \mem[2][15]~q ;
wire \mem[1][15]~q ;
wire \mem[7][47]~q ;
wire \mem~67_combout ;
wire \mem[6][47]~q ;
wire \mem[5][47]~q ;
wire \mem[4][47]~q ;
wire \mem[3][47]~q ;
wire \mem[2][47]~q ;
wire \mem[1][47]~q ;
wire \mem[7][23]~q ;
wire \mem~68_combout ;
wire \mem[6][23]~q ;
wire \mem[5][23]~q ;
wire \mem[4][23]~q ;
wire \mem[3][23]~q ;
wire \mem[2][23]~q ;
wire \mem[1][23]~q ;
wire \mem[7][55]~q ;
wire \mem~69_combout ;
wire \mem[6][55]~q ;
wire \mem[5][55]~q ;
wire \mem[4][55]~q ;
wire \mem[3][55]~q ;
wire \mem[2][55]~q ;
wire \mem[1][55]~q ;
wire \mem[7][31]~q ;
wire \mem~70_combout ;
wire \mem[6][31]~q ;
wire \mem[5][31]~q ;
wire \mem[4][31]~q ;
wire \mem[3][31]~q ;
wire \mem[2][31]~q ;
wire \mem[1][31]~q ;
wire \mem[7][63]~q ;
wire \mem~71_combout ;
wire \mem[6][63]~q ;
wire \mem[5][63]~q ;
wire \mem[4][63]~q ;
wire \mem[3][63]~q ;
wire \mem[2][63]~q ;
wire \mem[1][63]~q ;
wire \mem[7][7]~q ;
wire \mem~72_combout ;
wire \mem[6][7]~q ;
wire \mem[5][7]~q ;
wire \mem[4][7]~q ;
wire \mem[3][7]~q ;
wire \mem[2][7]~q ;
wire \mem[1][7]~q ;
wire \mem[7][39]~q ;
wire \mem~73_combout ;
wire \mem[6][39]~q ;
wire \mem[5][39]~q ;
wire \mem[4][39]~q ;
wire \mem[3][39]~q ;
wire \mem[2][39]~q ;
wire \mem[1][39]~q ;
wire \mem_used[7]~0_combout ;
wire \mem_used[0]~1_combout ;


dffeas \mem[0][105] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[1][105]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][139] (
	.clk(clk),
	.d(saved_grant_1),
	.asdata(\mem[1][139]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_139_0),
	.prn(vcc));
defparam \mem[0][139] .is_wysiwyg = "true";
defparam \mem[0][139] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(ShiftLeft04),
	.asdata(\mem[1][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[1][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_64_0),
	.prn(vcc));
defparam \mem[0][64] .is_wysiwyg = "true";
defparam \mem[0][64] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(ShiftLeft05),
	.asdata(\mem[1][69]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(ShiftLeft01),
	.asdata(\mem[1][65]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][70] (
	.clk(clk),
	.d(ShiftLeft06),
	.asdata(\mem[1][70]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_70_0),
	.prn(vcc));
defparam \mem[0][70] .is_wysiwyg = "true";
defparam \mem[0][70] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(ShiftLeft02),
	.asdata(\mem[1][66]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][71] (
	.clk(clk),
	.d(ShiftLeft07),
	.asdata(\mem[1][71]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_71_0),
	.prn(vcc));
defparam \mem[0][71] .is_wysiwyg = "true";
defparam \mem[0][71] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(ShiftLeft03),
	.asdata(\mem[1][67]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(ShiftLeft18),
	.asdata(\mem[1][8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][40] (
	.clk(clk),
	.d(ShiftLeft140),
	.asdata(\mem[1][40]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_40_0),
	.prn(vcc));
defparam \mem[0][40] .is_wysiwyg = "true";
defparam \mem[0][40] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(ShiftLeft116),
	.asdata(\mem[1][16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][48] (
	.clk(clk),
	.d(ShiftLeft148),
	.asdata(\mem[1][48]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_48_0),
	.prn(vcc));
defparam \mem[0][48] .is_wysiwyg = "true";
defparam \mem[0][48] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(ShiftLeft124),
	.asdata(\mem[1][24]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(ShiftLeft156),
	.asdata(\mem[1][56]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem[0][0] (
	.clk(clk),
	.d(ShiftLeft1),
	.asdata(\mem[1][0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][32] (
	.clk(clk),
	.d(ShiftLeft132),
	.asdata(\mem[1][32]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_32_0),
	.prn(vcc));
defparam \mem[0][32] .is_wysiwyg = "true";
defparam \mem[0][32] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(ShiftLeft19),
	.asdata(\mem[1][9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][41] (
	.clk(clk),
	.d(ShiftLeft141),
	.asdata(\mem[1][41]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_41_0),
	.prn(vcc));
defparam \mem[0][41] .is_wysiwyg = "true";
defparam \mem[0][41] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(ShiftLeft117),
	.asdata(\mem[1][17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][49] (
	.clk(clk),
	.d(ShiftLeft149),
	.asdata(\mem[1][49]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_49_0),
	.prn(vcc));
defparam \mem[0][49] .is_wysiwyg = "true";
defparam \mem[0][49] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(ShiftLeft125),
	.asdata(\mem[1][25]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(ShiftLeft157),
	.asdata(\mem[1][57]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(ShiftLeft11),
	.asdata(\mem[1][1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][33] (
	.clk(clk),
	.d(ShiftLeft133),
	.asdata(\mem[1][33]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_33_0),
	.prn(vcc));
defparam \mem[0][33] .is_wysiwyg = "true";
defparam \mem[0][33] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(ShiftLeft110),
	.asdata(\mem[1][10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][42] (
	.clk(clk),
	.d(ShiftLeft142),
	.asdata(\mem[1][42]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_42_0),
	.prn(vcc));
defparam \mem[0][42] .is_wysiwyg = "true";
defparam \mem[0][42] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(ShiftLeft118),
	.asdata(\mem[1][18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][50] (
	.clk(clk),
	.d(ShiftLeft150),
	.asdata(\mem[1][50]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_50_0),
	.prn(vcc));
defparam \mem[0][50] .is_wysiwyg = "true";
defparam \mem[0][50] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(ShiftLeft126),
	.asdata(\mem[1][26]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][58] (
	.clk(clk),
	.d(ShiftLeft158),
	.asdata(\mem[1][58]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_58_0),
	.prn(vcc));
defparam \mem[0][58] .is_wysiwyg = "true";
defparam \mem[0][58] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(ShiftLeft12),
	.asdata(\mem[1][2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][34] (
	.clk(clk),
	.d(ShiftLeft134),
	.asdata(\mem[1][34]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_34_0),
	.prn(vcc));
defparam \mem[0][34] .is_wysiwyg = "true";
defparam \mem[0][34] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(ShiftLeft111),
	.asdata(\mem[1][11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][43] (
	.clk(clk),
	.d(ShiftLeft143),
	.asdata(\mem[1][43]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_43_0),
	.prn(vcc));
defparam \mem[0][43] .is_wysiwyg = "true";
defparam \mem[0][43] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(ShiftLeft119),
	.asdata(\mem[1][19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][51] (
	.clk(clk),
	.d(ShiftLeft151),
	.asdata(\mem[1][51]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_51_0),
	.prn(vcc));
defparam \mem[0][51] .is_wysiwyg = "true";
defparam \mem[0][51] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(ShiftLeft127),
	.asdata(\mem[1][27]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(ShiftLeft159),
	.asdata(\mem[1][59]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(ShiftLeft13),
	.asdata(\mem[1][3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][35] (
	.clk(clk),
	.d(ShiftLeft135),
	.asdata(\mem[1][35]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_35_0),
	.prn(vcc));
defparam \mem[0][35] .is_wysiwyg = "true";
defparam \mem[0][35] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(ShiftLeft112),
	.asdata(\mem[1][12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][44] (
	.clk(clk),
	.d(ShiftLeft144),
	.asdata(\mem[1][44]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_44_0),
	.prn(vcc));
defparam \mem[0][44] .is_wysiwyg = "true";
defparam \mem[0][44] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(ShiftLeft120),
	.asdata(\mem[1][20]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][52] (
	.clk(clk),
	.d(ShiftLeft152),
	.asdata(\mem[1][52]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_52_0),
	.prn(vcc));
defparam \mem[0][52] .is_wysiwyg = "true";
defparam \mem[0][52] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(ShiftLeft128),
	.asdata(\mem[1][28]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][60] (
	.clk(clk),
	.d(ShiftLeft160),
	.asdata(\mem[1][60]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_60_0),
	.prn(vcc));
defparam \mem[0][60] .is_wysiwyg = "true";
defparam \mem[0][60] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(ShiftLeft14),
	.asdata(\mem[1][4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][36] (
	.clk(clk),
	.d(ShiftLeft136),
	.asdata(\mem[1][36]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_36_0),
	.prn(vcc));
defparam \mem[0][36] .is_wysiwyg = "true";
defparam \mem[0][36] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(ShiftLeft113),
	.asdata(\mem[1][13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][45] (
	.clk(clk),
	.d(ShiftLeft145),
	.asdata(\mem[1][45]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_45_0),
	.prn(vcc));
defparam \mem[0][45] .is_wysiwyg = "true";
defparam \mem[0][45] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(ShiftLeft121),
	.asdata(\mem[1][21]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][53] (
	.clk(clk),
	.d(ShiftLeft153),
	.asdata(\mem[1][53]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_53_0),
	.prn(vcc));
defparam \mem[0][53] .is_wysiwyg = "true";
defparam \mem[0][53] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(ShiftLeft129),
	.asdata(\mem[1][29]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(ShiftLeft161),
	.asdata(\mem[1][61]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(ShiftLeft15),
	.asdata(\mem[1][5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][37] (
	.clk(clk),
	.d(ShiftLeft137),
	.asdata(\mem[1][37]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_37_0),
	.prn(vcc));
defparam \mem[0][37] .is_wysiwyg = "true";
defparam \mem[0][37] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(ShiftLeft114),
	.asdata(\mem[1][14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][46] (
	.clk(clk),
	.d(ShiftLeft146),
	.asdata(\mem[1][46]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_46_0),
	.prn(vcc));
defparam \mem[0][46] .is_wysiwyg = "true";
defparam \mem[0][46] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(ShiftLeft122),
	.asdata(\mem[1][22]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][54] (
	.clk(clk),
	.d(ShiftLeft154),
	.asdata(\mem[1][54]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_54_0),
	.prn(vcc));
defparam \mem[0][54] .is_wysiwyg = "true";
defparam \mem[0][54] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(ShiftLeft130),
	.asdata(\mem[1][30]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][62] (
	.clk(clk),
	.d(ShiftLeft162),
	.asdata(\mem[1][62]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_62_0),
	.prn(vcc));
defparam \mem[0][62] .is_wysiwyg = "true";
defparam \mem[0][62] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(ShiftLeft16),
	.asdata(\mem[1][6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][38] (
	.clk(clk),
	.d(ShiftLeft138),
	.asdata(\mem[1][38]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_38_0),
	.prn(vcc));
defparam \mem[0][38] .is_wysiwyg = "true";
defparam \mem[0][38] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(ShiftLeft115),
	.asdata(\mem[1][15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][47] (
	.clk(clk),
	.d(ShiftLeft147),
	.asdata(\mem[1][47]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_47_0),
	.prn(vcc));
defparam \mem[0][47] .is_wysiwyg = "true";
defparam \mem[0][47] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(ShiftLeft123),
	.asdata(\mem[1][23]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][55] (
	.clk(clk),
	.d(ShiftLeft155),
	.asdata(\mem[1][55]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_55_0),
	.prn(vcc));
defparam \mem[0][55] .is_wysiwyg = "true";
defparam \mem[0][55] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(ShiftLeft131),
	.asdata(\mem[1][31]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

dffeas \mem[0][63] (
	.clk(clk),
	.d(ShiftLeft163),
	.asdata(\mem[1][63]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_63_0),
	.prn(vcc));
defparam \mem[0][63] .is_wysiwyg = "true";
defparam \mem[0][63] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(ShiftLeft17),
	.asdata(\mem[1][7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][39] (
	.clk(clk),
	.d(ShiftLeft139),
	.asdata(\mem[1][39]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[1]~q ),
	.ena(\always0~0_combout ),
	.q(mem_39_0),
	.prn(vcc));
defparam \mem[0][39] .is_wysiwyg = "true";
defparam \mem[0][39] .power_up = "low";

dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used[7]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_7),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[7][106] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][106]~q ),
	.prn(vcc));
defparam \mem[7][106] .is_wysiwyg = "true";
defparam \mem[7][106] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_7),
	.datab(!src_payload),
	.datac(!\mem[7][106]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_7),
	.datab(!src_valid),
	.datac(!write_cp_ready),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0202020202020202;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used~4 (
	.dataa(!mem_used_0),
	.datab(!\write~0_combout ),
	.datac(!\mem_used[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~4 .extended_lut = "off";
defparam \mem_used~4 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \mem_used~4 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[6]~3 (
	.dataa(!bready),
	.datab(!\write~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[6]~3 .extended_lut = "off";
defparam \mem_used[6]~3 .lut_mask = 64'h6666666666666666;
defparam \mem_used[6]~3 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used~6 (
	.dataa(!\write~0_combout ),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~6 .extended_lut = "off";
defparam \mem_used~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_used~6 .shared_arith = "off";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cyclonev_lcell_comb \mem_used~8 (
	.dataa(!\write~0_combout ),
	.datab(!\mem_used[2]~q ),
	.datac(!\mem_used[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~8 .extended_lut = "off";
defparam \mem_used~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_used~8 .shared_arith = "off";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cyclonev_lcell_comb \mem_used~7 (
	.dataa(!\write~0_combout ),
	.datab(!\mem_used[5]~q ),
	.datac(!\mem_used[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~7 .extended_lut = "off";
defparam \mem_used~7 .lut_mask = 64'h2727272727272727;
defparam \mem_used~7 .shared_arith = "off";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cyclonev_lcell_comb \mem_used~5 (
	.dataa(!\write~0_combout ),
	.datab(!\mem_used[6]~q ),
	.datac(!\mem_used[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~5 .extended_lut = "off";
defparam \mem_used~5 .lut_mask = 64'h2727272727272727;
defparam \mem_used~5 .shared_arith = "off";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cyclonev_lcell_comb \mem_used~2 (
	.dataa(!mem_used_7),
	.datab(!\write~0_combout ),
	.datac(!\mem_used[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used~2 .extended_lut = "off";
defparam \mem_used~2 .lut_mask = 64'h5757575757575757;
defparam \mem_used~2 .shared_arith = "off";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[6]~3_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cyclonev_lcell_comb \always6~0 (
	.dataa(!bready),
	.datab(!\mem_used[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always6~0 .shared_arith = "off";

dffeas \mem[6][105] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][105]~q ),
	.prn(vcc));
defparam \mem[6][105] .is_wysiwyg = "true";
defparam \mem[6][105] .power_up = "low";

cyclonev_lcell_comb \always5~0 (
	.dataa(!bready),
	.datab(!\mem_used[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always5~0 .shared_arith = "off";

dffeas \mem[5][105] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[6][105]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][105]~q ),
	.prn(vcc));
defparam \mem[5][105] .is_wysiwyg = "true";
defparam \mem[5][105] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!bready),
	.datab(!\mem_used[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[4][105] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[5][105]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][105]~q ),
	.prn(vcc));
defparam \mem[4][105] .is_wysiwyg = "true";
defparam \mem[4][105] .power_up = "low";

cyclonev_lcell_comb \always3~0 (
	.dataa(!bready),
	.datab(!\mem_used[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always3~0 .shared_arith = "off";

dffeas \mem[3][105] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[4][105]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][105]~q ),
	.prn(vcc));
defparam \mem[3][105] .is_wysiwyg = "true";
defparam \mem[3][105] .power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!bready),
	.datab(!\mem_used[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always2~0 .shared_arith = "off";

dffeas \mem[2][105] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[3][105]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][105]~q ),
	.prn(vcc));
defparam \mem[2][105] .is_wysiwyg = "true";
defparam \mem[2][105] .power_up = "low";

cyclonev_lcell_comb \always1~0 (
	.dataa(!bready),
	.datab(!\mem_used[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always1~0 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(src_payload),
	.asdata(\mem[2][105]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[7][154] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][154]~q ),
	.prn(vcc));
defparam \mem[7][154] .is_wysiwyg = "true";
defparam \mem[7][154] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_7),
	.datab(!saved_grant_1),
	.datac(!\mem[7][154]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[6][139] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][139]~q ),
	.prn(vcc));
defparam \mem[6][139] .is_wysiwyg = "true";
defparam \mem[6][139] .power_up = "low";

dffeas \mem[5][139] (
	.clk(clk),
	.d(saved_grant_1),
	.asdata(\mem[6][139]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][139]~q ),
	.prn(vcc));
defparam \mem[5][139] .is_wysiwyg = "true";
defparam \mem[5][139] .power_up = "low";

dffeas \mem[4][139] (
	.clk(clk),
	.d(saved_grant_1),
	.asdata(\mem[5][139]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][139]~q ),
	.prn(vcc));
defparam \mem[4][139] .is_wysiwyg = "true";
defparam \mem[4][139] .power_up = "low";

dffeas \mem[3][139] (
	.clk(clk),
	.d(saved_grant_1),
	.asdata(\mem[4][139]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][139]~q ),
	.prn(vcc));
defparam \mem[3][139] .is_wysiwyg = "true";
defparam \mem[3][139] .power_up = "low";

dffeas \mem[2][139] (
	.clk(clk),
	.d(saved_grant_1),
	.asdata(\mem[3][139]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][139]~q ),
	.prn(vcc));
defparam \mem[2][139] .is_wysiwyg = "true";
defparam \mem[2][139] .power_up = "low";

dffeas \mem[1][139] (
	.clk(clk),
	.d(saved_grant_1),
	.asdata(\mem[2][139]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][139]~q ),
	.prn(vcc));
defparam \mem[1][139] .is_wysiwyg = "true";
defparam \mem[1][139] .power_up = "low";

dffeas \mem[7][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][68]~q ),
	.prn(vcc));
defparam \mem[7][68] .is_wysiwyg = "true";
defparam \mem[7][68] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft04),
	.datac(!\mem[7][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[6][68] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][68]~q ),
	.prn(vcc));
defparam \mem[6][68] .is_wysiwyg = "true";
defparam \mem[6][68] .power_up = "low";

dffeas \mem[5][68] (
	.clk(clk),
	.d(ShiftLeft04),
	.asdata(\mem[6][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][68]~q ),
	.prn(vcc));
defparam \mem[5][68] .is_wysiwyg = "true";
defparam \mem[5][68] .power_up = "low";

dffeas \mem[4][68] (
	.clk(clk),
	.d(ShiftLeft04),
	.asdata(\mem[5][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][68]~q ),
	.prn(vcc));
defparam \mem[4][68] .is_wysiwyg = "true";
defparam \mem[4][68] .power_up = "low";

dffeas \mem[3][68] (
	.clk(clk),
	.d(ShiftLeft04),
	.asdata(\mem[4][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][68]~q ),
	.prn(vcc));
defparam \mem[3][68] .is_wysiwyg = "true";
defparam \mem[3][68] .power_up = "low";

dffeas \mem[2][68] (
	.clk(clk),
	.d(ShiftLeft04),
	.asdata(\mem[3][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][68]~q ),
	.prn(vcc));
defparam \mem[2][68] .is_wysiwyg = "true";
defparam \mem[2][68] .power_up = "low";

dffeas \mem[1][68] (
	.clk(clk),
	.d(ShiftLeft04),
	.asdata(\mem[2][68]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

dffeas \mem[7][64] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][64]~q ),
	.prn(vcc));
defparam \mem[7][64] .is_wysiwyg = "true";
defparam \mem[7][64] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft0),
	.datac(!\mem[7][64]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h2727272727272727;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[6][64] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][64]~q ),
	.prn(vcc));
defparam \mem[6][64] .is_wysiwyg = "true";
defparam \mem[6][64] .power_up = "low";

dffeas \mem[5][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[6][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][64]~q ),
	.prn(vcc));
defparam \mem[5][64] .is_wysiwyg = "true";
defparam \mem[5][64] .power_up = "low";

dffeas \mem[4][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[5][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][64]~q ),
	.prn(vcc));
defparam \mem[4][64] .is_wysiwyg = "true";
defparam \mem[4][64] .power_up = "low";

dffeas \mem[3][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[4][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][64]~q ),
	.prn(vcc));
defparam \mem[3][64] .is_wysiwyg = "true";
defparam \mem[3][64] .power_up = "low";

dffeas \mem[2][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[3][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][64]~q ),
	.prn(vcc));
defparam \mem[2][64] .is_wysiwyg = "true";
defparam \mem[2][64] .power_up = "low";

dffeas \mem[1][64] (
	.clk(clk),
	.d(ShiftLeft0),
	.asdata(\mem[2][64]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][64]~q ),
	.prn(vcc));
defparam \mem[1][64] .is_wysiwyg = "true";
defparam \mem[1][64] .power_up = "low";

dffeas \mem[7][69] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][69]~q ),
	.prn(vcc));
defparam \mem[7][69] .is_wysiwyg = "true";
defparam \mem[7][69] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft05),
	.datac(!\mem[7][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h2727272727272727;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[6][69] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][69]~q ),
	.prn(vcc));
defparam \mem[6][69] .is_wysiwyg = "true";
defparam \mem[6][69] .power_up = "low";

dffeas \mem[5][69] (
	.clk(clk),
	.d(ShiftLeft05),
	.asdata(\mem[6][69]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][69]~q ),
	.prn(vcc));
defparam \mem[5][69] .is_wysiwyg = "true";
defparam \mem[5][69] .power_up = "low";

dffeas \mem[4][69] (
	.clk(clk),
	.d(ShiftLeft05),
	.asdata(\mem[5][69]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][69]~q ),
	.prn(vcc));
defparam \mem[4][69] .is_wysiwyg = "true";
defparam \mem[4][69] .power_up = "low";

dffeas \mem[3][69] (
	.clk(clk),
	.d(ShiftLeft05),
	.asdata(\mem[4][69]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][69]~q ),
	.prn(vcc));
defparam \mem[3][69] .is_wysiwyg = "true";
defparam \mem[3][69] .power_up = "low";

dffeas \mem[2][69] (
	.clk(clk),
	.d(ShiftLeft05),
	.asdata(\mem[3][69]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][69]~q ),
	.prn(vcc));
defparam \mem[2][69] .is_wysiwyg = "true";
defparam \mem[2][69] .power_up = "low";

dffeas \mem[1][69] (
	.clk(clk),
	.d(ShiftLeft05),
	.asdata(\mem[2][69]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

dffeas \mem[7][65] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][65]~q ),
	.prn(vcc));
defparam \mem[7][65] .is_wysiwyg = "true";
defparam \mem[7][65] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft01),
	.datac(!\mem[7][65]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h2727272727272727;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[6][65] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][65]~q ),
	.prn(vcc));
defparam \mem[6][65] .is_wysiwyg = "true";
defparam \mem[6][65] .power_up = "low";

dffeas \mem[5][65] (
	.clk(clk),
	.d(ShiftLeft01),
	.asdata(\mem[6][65]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][65]~q ),
	.prn(vcc));
defparam \mem[5][65] .is_wysiwyg = "true";
defparam \mem[5][65] .power_up = "low";

dffeas \mem[4][65] (
	.clk(clk),
	.d(ShiftLeft01),
	.asdata(\mem[5][65]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][65]~q ),
	.prn(vcc));
defparam \mem[4][65] .is_wysiwyg = "true";
defparam \mem[4][65] .power_up = "low";

dffeas \mem[3][65] (
	.clk(clk),
	.d(ShiftLeft01),
	.asdata(\mem[4][65]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][65]~q ),
	.prn(vcc));
defparam \mem[3][65] .is_wysiwyg = "true";
defparam \mem[3][65] .power_up = "low";

dffeas \mem[2][65] (
	.clk(clk),
	.d(ShiftLeft01),
	.asdata(\mem[3][65]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][65]~q ),
	.prn(vcc));
defparam \mem[2][65] .is_wysiwyg = "true";
defparam \mem[2][65] .power_up = "low";

dffeas \mem[1][65] (
	.clk(clk),
	.d(ShiftLeft01),
	.asdata(\mem[2][65]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

dffeas \mem[7][70] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][70]~q ),
	.prn(vcc));
defparam \mem[7][70] .is_wysiwyg = "true";
defparam \mem[7][70] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft06),
	.datac(!\mem[7][70]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h2727272727272727;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[6][70] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][70]~q ),
	.prn(vcc));
defparam \mem[6][70] .is_wysiwyg = "true";
defparam \mem[6][70] .power_up = "low";

dffeas \mem[5][70] (
	.clk(clk),
	.d(ShiftLeft06),
	.asdata(\mem[6][70]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][70]~q ),
	.prn(vcc));
defparam \mem[5][70] .is_wysiwyg = "true";
defparam \mem[5][70] .power_up = "low";

dffeas \mem[4][70] (
	.clk(clk),
	.d(ShiftLeft06),
	.asdata(\mem[5][70]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][70]~q ),
	.prn(vcc));
defparam \mem[4][70] .is_wysiwyg = "true";
defparam \mem[4][70] .power_up = "low";

dffeas \mem[3][70] (
	.clk(clk),
	.d(ShiftLeft06),
	.asdata(\mem[4][70]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][70]~q ),
	.prn(vcc));
defparam \mem[3][70] .is_wysiwyg = "true";
defparam \mem[3][70] .power_up = "low";

dffeas \mem[2][70] (
	.clk(clk),
	.d(ShiftLeft06),
	.asdata(\mem[3][70]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][70]~q ),
	.prn(vcc));
defparam \mem[2][70] .is_wysiwyg = "true";
defparam \mem[2][70] .power_up = "low";

dffeas \mem[1][70] (
	.clk(clk),
	.d(ShiftLeft06),
	.asdata(\mem[2][70]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][70]~q ),
	.prn(vcc));
defparam \mem[1][70] .is_wysiwyg = "true";
defparam \mem[1][70] .power_up = "low";

dffeas \mem[7][66] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][66]~q ),
	.prn(vcc));
defparam \mem[7][66] .is_wysiwyg = "true";
defparam \mem[7][66] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft02),
	.datac(!\mem[7][66]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h2727272727272727;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[6][66] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][66]~q ),
	.prn(vcc));
defparam \mem[6][66] .is_wysiwyg = "true";
defparam \mem[6][66] .power_up = "low";

dffeas \mem[5][66] (
	.clk(clk),
	.d(ShiftLeft02),
	.asdata(\mem[6][66]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][66]~q ),
	.prn(vcc));
defparam \mem[5][66] .is_wysiwyg = "true";
defparam \mem[5][66] .power_up = "low";

dffeas \mem[4][66] (
	.clk(clk),
	.d(ShiftLeft02),
	.asdata(\mem[5][66]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][66]~q ),
	.prn(vcc));
defparam \mem[4][66] .is_wysiwyg = "true";
defparam \mem[4][66] .power_up = "low";

dffeas \mem[3][66] (
	.clk(clk),
	.d(ShiftLeft02),
	.asdata(\mem[4][66]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][66]~q ),
	.prn(vcc));
defparam \mem[3][66] .is_wysiwyg = "true";
defparam \mem[3][66] .power_up = "low";

dffeas \mem[2][66] (
	.clk(clk),
	.d(ShiftLeft02),
	.asdata(\mem[3][66]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][66]~q ),
	.prn(vcc));
defparam \mem[2][66] .is_wysiwyg = "true";
defparam \mem[2][66] .power_up = "low";

dffeas \mem[1][66] (
	.clk(clk),
	.d(ShiftLeft02),
	.asdata(\mem[2][66]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

dffeas \mem[7][71] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][71]~q ),
	.prn(vcc));
defparam \mem[7][71] .is_wysiwyg = "true";
defparam \mem[7][71] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft07),
	.datac(!\mem[7][71]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h2727272727272727;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[6][71] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][71]~q ),
	.prn(vcc));
defparam \mem[6][71] .is_wysiwyg = "true";
defparam \mem[6][71] .power_up = "low";

dffeas \mem[5][71] (
	.clk(clk),
	.d(ShiftLeft07),
	.asdata(\mem[6][71]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][71]~q ),
	.prn(vcc));
defparam \mem[5][71] .is_wysiwyg = "true";
defparam \mem[5][71] .power_up = "low";

dffeas \mem[4][71] (
	.clk(clk),
	.d(ShiftLeft07),
	.asdata(\mem[5][71]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][71]~q ),
	.prn(vcc));
defparam \mem[4][71] .is_wysiwyg = "true";
defparam \mem[4][71] .power_up = "low";

dffeas \mem[3][71] (
	.clk(clk),
	.d(ShiftLeft07),
	.asdata(\mem[4][71]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][71]~q ),
	.prn(vcc));
defparam \mem[3][71] .is_wysiwyg = "true";
defparam \mem[3][71] .power_up = "low";

dffeas \mem[2][71] (
	.clk(clk),
	.d(ShiftLeft07),
	.asdata(\mem[3][71]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][71]~q ),
	.prn(vcc));
defparam \mem[2][71] .is_wysiwyg = "true";
defparam \mem[2][71] .power_up = "low";

dffeas \mem[1][71] (
	.clk(clk),
	.d(ShiftLeft07),
	.asdata(\mem[2][71]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][71]~q ),
	.prn(vcc));
defparam \mem[1][71] .is_wysiwyg = "true";
defparam \mem[1][71] .power_up = "low";

dffeas \mem[7][67] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][67]~q ),
	.prn(vcc));
defparam \mem[7][67] .is_wysiwyg = "true";
defparam \mem[7][67] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft03),
	.datac(!\mem[7][67]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h2727272727272727;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[6][67] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][67]~q ),
	.prn(vcc));
defparam \mem[6][67] .is_wysiwyg = "true";
defparam \mem[6][67] .power_up = "low";

dffeas \mem[5][67] (
	.clk(clk),
	.d(ShiftLeft03),
	.asdata(\mem[6][67]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][67]~q ),
	.prn(vcc));
defparam \mem[5][67] .is_wysiwyg = "true";
defparam \mem[5][67] .power_up = "low";

dffeas \mem[4][67] (
	.clk(clk),
	.d(ShiftLeft03),
	.asdata(\mem[5][67]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][67]~q ),
	.prn(vcc));
defparam \mem[4][67] .is_wysiwyg = "true";
defparam \mem[4][67] .power_up = "low";

dffeas \mem[3][67] (
	.clk(clk),
	.d(ShiftLeft03),
	.asdata(\mem[4][67]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][67]~q ),
	.prn(vcc));
defparam \mem[3][67] .is_wysiwyg = "true";
defparam \mem[3][67] .power_up = "low";

dffeas \mem[2][67] (
	.clk(clk),
	.d(ShiftLeft03),
	.asdata(\mem[3][67]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][67]~q ),
	.prn(vcc));
defparam \mem[2][67] .is_wysiwyg = "true";
defparam \mem[2][67] .power_up = "low";

dffeas \mem[1][67] (
	.clk(clk),
	.d(ShiftLeft03),
	.asdata(\mem[2][67]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

dffeas \mem[7][8] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][8]~q ),
	.prn(vcc));
defparam \mem[7][8] .is_wysiwyg = "true";
defparam \mem[7][8] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft18),
	.datac(!\mem[7][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h2727272727272727;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[6][8] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][8]~q ),
	.prn(vcc));
defparam \mem[6][8] .is_wysiwyg = "true";
defparam \mem[6][8] .power_up = "low";

dffeas \mem[5][8] (
	.clk(clk),
	.d(ShiftLeft18),
	.asdata(\mem[6][8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][8]~q ),
	.prn(vcc));
defparam \mem[5][8] .is_wysiwyg = "true";
defparam \mem[5][8] .power_up = "low";

dffeas \mem[4][8] (
	.clk(clk),
	.d(ShiftLeft18),
	.asdata(\mem[5][8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][8]~q ),
	.prn(vcc));
defparam \mem[4][8] .is_wysiwyg = "true";
defparam \mem[4][8] .power_up = "low";

dffeas \mem[3][8] (
	.clk(clk),
	.d(ShiftLeft18),
	.asdata(\mem[4][8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][8]~q ),
	.prn(vcc));
defparam \mem[3][8] .is_wysiwyg = "true";
defparam \mem[3][8] .power_up = "low";

dffeas \mem[2][8] (
	.clk(clk),
	.d(ShiftLeft18),
	.asdata(\mem[3][8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][8]~q ),
	.prn(vcc));
defparam \mem[2][8] .is_wysiwyg = "true";
defparam \mem[2][8] .power_up = "low";

dffeas \mem[1][8] (
	.clk(clk),
	.d(ShiftLeft18),
	.asdata(\mem[2][8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

dffeas \mem[7][40] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][40]~q ),
	.prn(vcc));
defparam \mem[7][40] .is_wysiwyg = "true";
defparam \mem[7][40] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft140),
	.datac(!\mem[7][40]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h2727272727272727;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[6][40] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][40]~q ),
	.prn(vcc));
defparam \mem[6][40] .is_wysiwyg = "true";
defparam \mem[6][40] .power_up = "low";

dffeas \mem[5][40] (
	.clk(clk),
	.d(ShiftLeft140),
	.asdata(\mem[6][40]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][40]~q ),
	.prn(vcc));
defparam \mem[5][40] .is_wysiwyg = "true";
defparam \mem[5][40] .power_up = "low";

dffeas \mem[4][40] (
	.clk(clk),
	.d(ShiftLeft140),
	.asdata(\mem[5][40]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][40]~q ),
	.prn(vcc));
defparam \mem[4][40] .is_wysiwyg = "true";
defparam \mem[4][40] .power_up = "low";

dffeas \mem[3][40] (
	.clk(clk),
	.d(ShiftLeft140),
	.asdata(\mem[4][40]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][40]~q ),
	.prn(vcc));
defparam \mem[3][40] .is_wysiwyg = "true";
defparam \mem[3][40] .power_up = "low";

dffeas \mem[2][40] (
	.clk(clk),
	.d(ShiftLeft140),
	.asdata(\mem[3][40]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][40]~q ),
	.prn(vcc));
defparam \mem[2][40] .is_wysiwyg = "true";
defparam \mem[2][40] .power_up = "low";

dffeas \mem[1][40] (
	.clk(clk),
	.d(ShiftLeft140),
	.asdata(\mem[2][40]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][40]~q ),
	.prn(vcc));
defparam \mem[1][40] .is_wysiwyg = "true";
defparam \mem[1][40] .power_up = "low";

dffeas \mem[7][16] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][16]~q ),
	.prn(vcc));
defparam \mem[7][16] .is_wysiwyg = "true";
defparam \mem[7][16] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft116),
	.datac(!\mem[7][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h2727272727272727;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[6][16] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][16]~q ),
	.prn(vcc));
defparam \mem[6][16] .is_wysiwyg = "true";
defparam \mem[6][16] .power_up = "low";

dffeas \mem[5][16] (
	.clk(clk),
	.d(ShiftLeft116),
	.asdata(\mem[6][16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][16]~q ),
	.prn(vcc));
defparam \mem[5][16] .is_wysiwyg = "true";
defparam \mem[5][16] .power_up = "low";

dffeas \mem[4][16] (
	.clk(clk),
	.d(ShiftLeft116),
	.asdata(\mem[5][16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][16]~q ),
	.prn(vcc));
defparam \mem[4][16] .is_wysiwyg = "true";
defparam \mem[4][16] .power_up = "low";

dffeas \mem[3][16] (
	.clk(clk),
	.d(ShiftLeft116),
	.asdata(\mem[4][16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][16]~q ),
	.prn(vcc));
defparam \mem[3][16] .is_wysiwyg = "true";
defparam \mem[3][16] .power_up = "low";

dffeas \mem[2][16] (
	.clk(clk),
	.d(ShiftLeft116),
	.asdata(\mem[3][16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][16]~q ),
	.prn(vcc));
defparam \mem[2][16] .is_wysiwyg = "true";
defparam \mem[2][16] .power_up = "low";

dffeas \mem[1][16] (
	.clk(clk),
	.d(ShiftLeft116),
	.asdata(\mem[2][16]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

dffeas \mem[7][48] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][48]~q ),
	.prn(vcc));
defparam \mem[7][48] .is_wysiwyg = "true";
defparam \mem[7][48] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft148),
	.datac(!\mem[7][48]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h2727272727272727;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[6][48] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][48]~q ),
	.prn(vcc));
defparam \mem[6][48] .is_wysiwyg = "true";
defparam \mem[6][48] .power_up = "low";

dffeas \mem[5][48] (
	.clk(clk),
	.d(ShiftLeft148),
	.asdata(\mem[6][48]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][48]~q ),
	.prn(vcc));
defparam \mem[5][48] .is_wysiwyg = "true";
defparam \mem[5][48] .power_up = "low";

dffeas \mem[4][48] (
	.clk(clk),
	.d(ShiftLeft148),
	.asdata(\mem[5][48]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][48]~q ),
	.prn(vcc));
defparam \mem[4][48] .is_wysiwyg = "true";
defparam \mem[4][48] .power_up = "low";

dffeas \mem[3][48] (
	.clk(clk),
	.d(ShiftLeft148),
	.asdata(\mem[4][48]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][48]~q ),
	.prn(vcc));
defparam \mem[3][48] .is_wysiwyg = "true";
defparam \mem[3][48] .power_up = "low";

dffeas \mem[2][48] (
	.clk(clk),
	.d(ShiftLeft148),
	.asdata(\mem[3][48]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][48]~q ),
	.prn(vcc));
defparam \mem[2][48] .is_wysiwyg = "true";
defparam \mem[2][48] .power_up = "low";

dffeas \mem[1][48] (
	.clk(clk),
	.d(ShiftLeft148),
	.asdata(\mem[2][48]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][48]~q ),
	.prn(vcc));
defparam \mem[1][48] .is_wysiwyg = "true";
defparam \mem[1][48] .power_up = "low";

dffeas \mem[7][24] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][24]~q ),
	.prn(vcc));
defparam \mem[7][24] .is_wysiwyg = "true";
defparam \mem[7][24] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft124),
	.datac(!\mem[7][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h2727272727272727;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[6][24] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][24]~q ),
	.prn(vcc));
defparam \mem[6][24] .is_wysiwyg = "true";
defparam \mem[6][24] .power_up = "low";

dffeas \mem[5][24] (
	.clk(clk),
	.d(ShiftLeft124),
	.asdata(\mem[6][24]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][24]~q ),
	.prn(vcc));
defparam \mem[5][24] .is_wysiwyg = "true";
defparam \mem[5][24] .power_up = "low";

dffeas \mem[4][24] (
	.clk(clk),
	.d(ShiftLeft124),
	.asdata(\mem[5][24]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][24]~q ),
	.prn(vcc));
defparam \mem[4][24] .is_wysiwyg = "true";
defparam \mem[4][24] .power_up = "low";

dffeas \mem[3][24] (
	.clk(clk),
	.d(ShiftLeft124),
	.asdata(\mem[4][24]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][24]~q ),
	.prn(vcc));
defparam \mem[3][24] .is_wysiwyg = "true";
defparam \mem[3][24] .power_up = "low";

dffeas \mem[2][24] (
	.clk(clk),
	.d(ShiftLeft124),
	.asdata(\mem[3][24]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][24]~q ),
	.prn(vcc));
defparam \mem[2][24] .is_wysiwyg = "true";
defparam \mem[2][24] .power_up = "low";

dffeas \mem[1][24] (
	.clk(clk),
	.d(ShiftLeft124),
	.asdata(\mem[2][24]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

dffeas \mem[7][56] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][56]~q ),
	.prn(vcc));
defparam \mem[7][56] .is_wysiwyg = "true";
defparam \mem[7][56] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft156),
	.datac(!\mem[7][56]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h2727272727272727;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[6][56] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][56]~q ),
	.prn(vcc));
defparam \mem[6][56] .is_wysiwyg = "true";
defparam \mem[6][56] .power_up = "low";

dffeas \mem[5][56] (
	.clk(clk),
	.d(ShiftLeft156),
	.asdata(\mem[6][56]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][56]~q ),
	.prn(vcc));
defparam \mem[5][56] .is_wysiwyg = "true";
defparam \mem[5][56] .power_up = "low";

dffeas \mem[4][56] (
	.clk(clk),
	.d(ShiftLeft156),
	.asdata(\mem[5][56]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][56]~q ),
	.prn(vcc));
defparam \mem[4][56] .is_wysiwyg = "true";
defparam \mem[4][56] .power_up = "low";

dffeas \mem[3][56] (
	.clk(clk),
	.d(ShiftLeft156),
	.asdata(\mem[4][56]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][56]~q ),
	.prn(vcc));
defparam \mem[3][56] .is_wysiwyg = "true";
defparam \mem[3][56] .power_up = "low";

dffeas \mem[2][56] (
	.clk(clk),
	.d(ShiftLeft156),
	.asdata(\mem[3][56]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][56]~q ),
	.prn(vcc));
defparam \mem[2][56] .is_wysiwyg = "true";
defparam \mem[2][56] .power_up = "low";

dffeas \mem[1][56] (
	.clk(clk),
	.d(ShiftLeft156),
	.asdata(\mem[2][56]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

dffeas \mem[7][0] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][0]~q ),
	.prn(vcc));
defparam \mem[7][0] .is_wysiwyg = "true";
defparam \mem[7][0] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft1),
	.datac(!\mem[7][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h2727272727272727;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[6][0] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][0]~q ),
	.prn(vcc));
defparam \mem[6][0] .is_wysiwyg = "true";
defparam \mem[6][0] .power_up = "low";

dffeas \mem[5][0] (
	.clk(clk),
	.d(ShiftLeft1),
	.asdata(\mem[6][0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][0]~q ),
	.prn(vcc));
defparam \mem[5][0] .is_wysiwyg = "true";
defparam \mem[5][0] .power_up = "low";

dffeas \mem[4][0] (
	.clk(clk),
	.d(ShiftLeft1),
	.asdata(\mem[5][0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][0]~q ),
	.prn(vcc));
defparam \mem[4][0] .is_wysiwyg = "true";
defparam \mem[4][0] .power_up = "low";

dffeas \mem[3][0] (
	.clk(clk),
	.d(ShiftLeft1),
	.asdata(\mem[4][0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][0]~q ),
	.prn(vcc));
defparam \mem[3][0] .is_wysiwyg = "true";
defparam \mem[3][0] .power_up = "low";

dffeas \mem[2][0] (
	.clk(clk),
	.d(ShiftLeft1),
	.asdata(\mem[3][0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][0]~q ),
	.prn(vcc));
defparam \mem[2][0] .is_wysiwyg = "true";
defparam \mem[2][0] .power_up = "low";

dffeas \mem[1][0] (
	.clk(clk),
	.d(ShiftLeft1),
	.asdata(\mem[2][0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

dffeas \mem[7][32] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][32]~q ),
	.prn(vcc));
defparam \mem[7][32] .is_wysiwyg = "true";
defparam \mem[7][32] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft132),
	.datac(!\mem[7][32]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h2727272727272727;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[6][32] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][32]~q ),
	.prn(vcc));
defparam \mem[6][32] .is_wysiwyg = "true";
defparam \mem[6][32] .power_up = "low";

dffeas \mem[5][32] (
	.clk(clk),
	.d(ShiftLeft132),
	.asdata(\mem[6][32]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][32]~q ),
	.prn(vcc));
defparam \mem[5][32] .is_wysiwyg = "true";
defparam \mem[5][32] .power_up = "low";

dffeas \mem[4][32] (
	.clk(clk),
	.d(ShiftLeft132),
	.asdata(\mem[5][32]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][32]~q ),
	.prn(vcc));
defparam \mem[4][32] .is_wysiwyg = "true";
defparam \mem[4][32] .power_up = "low";

dffeas \mem[3][32] (
	.clk(clk),
	.d(ShiftLeft132),
	.asdata(\mem[4][32]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][32]~q ),
	.prn(vcc));
defparam \mem[3][32] .is_wysiwyg = "true";
defparam \mem[3][32] .power_up = "low";

dffeas \mem[2][32] (
	.clk(clk),
	.d(ShiftLeft132),
	.asdata(\mem[3][32]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][32]~q ),
	.prn(vcc));
defparam \mem[2][32] .is_wysiwyg = "true";
defparam \mem[2][32] .power_up = "low";

dffeas \mem[1][32] (
	.clk(clk),
	.d(ShiftLeft132),
	.asdata(\mem[2][32]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][32]~q ),
	.prn(vcc));
defparam \mem[1][32] .is_wysiwyg = "true";
defparam \mem[1][32] .power_up = "low";

dffeas \mem[7][9] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][9]~q ),
	.prn(vcc));
defparam \mem[7][9] .is_wysiwyg = "true";
defparam \mem[7][9] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft19),
	.datac(!\mem[7][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h2727272727272727;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[6][9] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][9]~q ),
	.prn(vcc));
defparam \mem[6][9] .is_wysiwyg = "true";
defparam \mem[6][9] .power_up = "low";

dffeas \mem[5][9] (
	.clk(clk),
	.d(ShiftLeft19),
	.asdata(\mem[6][9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][9]~q ),
	.prn(vcc));
defparam \mem[5][9] .is_wysiwyg = "true";
defparam \mem[5][9] .power_up = "low";

dffeas \mem[4][9] (
	.clk(clk),
	.d(ShiftLeft19),
	.asdata(\mem[5][9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][9]~q ),
	.prn(vcc));
defparam \mem[4][9] .is_wysiwyg = "true";
defparam \mem[4][9] .power_up = "low";

dffeas \mem[3][9] (
	.clk(clk),
	.d(ShiftLeft19),
	.asdata(\mem[4][9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][9]~q ),
	.prn(vcc));
defparam \mem[3][9] .is_wysiwyg = "true";
defparam \mem[3][9] .power_up = "low";

dffeas \mem[2][9] (
	.clk(clk),
	.d(ShiftLeft19),
	.asdata(\mem[3][9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][9]~q ),
	.prn(vcc));
defparam \mem[2][9] .is_wysiwyg = "true";
defparam \mem[2][9] .power_up = "low";

dffeas \mem[1][9] (
	.clk(clk),
	.d(ShiftLeft19),
	.asdata(\mem[2][9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

dffeas \mem[7][41] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][41]~q ),
	.prn(vcc));
defparam \mem[7][41] .is_wysiwyg = "true";
defparam \mem[7][41] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft141),
	.datac(!\mem[7][41]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h2727272727272727;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[6][41] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][41]~q ),
	.prn(vcc));
defparam \mem[6][41] .is_wysiwyg = "true";
defparam \mem[6][41] .power_up = "low";

dffeas \mem[5][41] (
	.clk(clk),
	.d(ShiftLeft141),
	.asdata(\mem[6][41]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][41]~q ),
	.prn(vcc));
defparam \mem[5][41] .is_wysiwyg = "true";
defparam \mem[5][41] .power_up = "low";

dffeas \mem[4][41] (
	.clk(clk),
	.d(ShiftLeft141),
	.asdata(\mem[5][41]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][41]~q ),
	.prn(vcc));
defparam \mem[4][41] .is_wysiwyg = "true";
defparam \mem[4][41] .power_up = "low";

dffeas \mem[3][41] (
	.clk(clk),
	.d(ShiftLeft141),
	.asdata(\mem[4][41]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][41]~q ),
	.prn(vcc));
defparam \mem[3][41] .is_wysiwyg = "true";
defparam \mem[3][41] .power_up = "low";

dffeas \mem[2][41] (
	.clk(clk),
	.d(ShiftLeft141),
	.asdata(\mem[3][41]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][41]~q ),
	.prn(vcc));
defparam \mem[2][41] .is_wysiwyg = "true";
defparam \mem[2][41] .power_up = "low";

dffeas \mem[1][41] (
	.clk(clk),
	.d(ShiftLeft141),
	.asdata(\mem[2][41]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][41]~q ),
	.prn(vcc));
defparam \mem[1][41] .is_wysiwyg = "true";
defparam \mem[1][41] .power_up = "low";

dffeas \mem[7][17] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][17]~q ),
	.prn(vcc));
defparam \mem[7][17] .is_wysiwyg = "true";
defparam \mem[7][17] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft117),
	.datac(!\mem[7][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h2727272727272727;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[6][17] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][17]~q ),
	.prn(vcc));
defparam \mem[6][17] .is_wysiwyg = "true";
defparam \mem[6][17] .power_up = "low";

dffeas \mem[5][17] (
	.clk(clk),
	.d(ShiftLeft117),
	.asdata(\mem[6][17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][17]~q ),
	.prn(vcc));
defparam \mem[5][17] .is_wysiwyg = "true";
defparam \mem[5][17] .power_up = "low";

dffeas \mem[4][17] (
	.clk(clk),
	.d(ShiftLeft117),
	.asdata(\mem[5][17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][17]~q ),
	.prn(vcc));
defparam \mem[4][17] .is_wysiwyg = "true";
defparam \mem[4][17] .power_up = "low";

dffeas \mem[3][17] (
	.clk(clk),
	.d(ShiftLeft117),
	.asdata(\mem[4][17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][17]~q ),
	.prn(vcc));
defparam \mem[3][17] .is_wysiwyg = "true";
defparam \mem[3][17] .power_up = "low";

dffeas \mem[2][17] (
	.clk(clk),
	.d(ShiftLeft117),
	.asdata(\mem[3][17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][17]~q ),
	.prn(vcc));
defparam \mem[2][17] .is_wysiwyg = "true";
defparam \mem[2][17] .power_up = "low";

dffeas \mem[1][17] (
	.clk(clk),
	.d(ShiftLeft117),
	.asdata(\mem[2][17]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

dffeas \mem[7][49] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][49]~q ),
	.prn(vcc));
defparam \mem[7][49] .is_wysiwyg = "true";
defparam \mem[7][49] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft149),
	.datac(!\mem[7][49]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h2727272727272727;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[6][49] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][49]~q ),
	.prn(vcc));
defparam \mem[6][49] .is_wysiwyg = "true";
defparam \mem[6][49] .power_up = "low";

dffeas \mem[5][49] (
	.clk(clk),
	.d(ShiftLeft149),
	.asdata(\mem[6][49]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][49]~q ),
	.prn(vcc));
defparam \mem[5][49] .is_wysiwyg = "true";
defparam \mem[5][49] .power_up = "low";

dffeas \mem[4][49] (
	.clk(clk),
	.d(ShiftLeft149),
	.asdata(\mem[5][49]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][49]~q ),
	.prn(vcc));
defparam \mem[4][49] .is_wysiwyg = "true";
defparam \mem[4][49] .power_up = "low";

dffeas \mem[3][49] (
	.clk(clk),
	.d(ShiftLeft149),
	.asdata(\mem[4][49]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][49]~q ),
	.prn(vcc));
defparam \mem[3][49] .is_wysiwyg = "true";
defparam \mem[3][49] .power_up = "low";

dffeas \mem[2][49] (
	.clk(clk),
	.d(ShiftLeft149),
	.asdata(\mem[3][49]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][49]~q ),
	.prn(vcc));
defparam \mem[2][49] .is_wysiwyg = "true";
defparam \mem[2][49] .power_up = "low";

dffeas \mem[1][49] (
	.clk(clk),
	.d(ShiftLeft149),
	.asdata(\mem[2][49]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][49]~q ),
	.prn(vcc));
defparam \mem[1][49] .is_wysiwyg = "true";
defparam \mem[1][49] .power_up = "low";

dffeas \mem[7][25] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][25]~q ),
	.prn(vcc));
defparam \mem[7][25] .is_wysiwyg = "true";
defparam \mem[7][25] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft125),
	.datac(!\mem[7][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h2727272727272727;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[6][25] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][25]~q ),
	.prn(vcc));
defparam \mem[6][25] .is_wysiwyg = "true";
defparam \mem[6][25] .power_up = "low";

dffeas \mem[5][25] (
	.clk(clk),
	.d(ShiftLeft125),
	.asdata(\mem[6][25]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][25]~q ),
	.prn(vcc));
defparam \mem[5][25] .is_wysiwyg = "true";
defparam \mem[5][25] .power_up = "low";

dffeas \mem[4][25] (
	.clk(clk),
	.d(ShiftLeft125),
	.asdata(\mem[5][25]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][25]~q ),
	.prn(vcc));
defparam \mem[4][25] .is_wysiwyg = "true";
defparam \mem[4][25] .power_up = "low";

dffeas \mem[3][25] (
	.clk(clk),
	.d(ShiftLeft125),
	.asdata(\mem[4][25]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][25]~q ),
	.prn(vcc));
defparam \mem[3][25] .is_wysiwyg = "true";
defparam \mem[3][25] .power_up = "low";

dffeas \mem[2][25] (
	.clk(clk),
	.d(ShiftLeft125),
	.asdata(\mem[3][25]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][25]~q ),
	.prn(vcc));
defparam \mem[2][25] .is_wysiwyg = "true";
defparam \mem[2][25] .power_up = "low";

dffeas \mem[1][25] (
	.clk(clk),
	.d(ShiftLeft125),
	.asdata(\mem[2][25]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

dffeas \mem[7][57] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][57]~q ),
	.prn(vcc));
defparam \mem[7][57] .is_wysiwyg = "true";
defparam \mem[7][57] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft157),
	.datac(!\mem[7][57]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h2727272727272727;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[6][57] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][57]~q ),
	.prn(vcc));
defparam \mem[6][57] .is_wysiwyg = "true";
defparam \mem[6][57] .power_up = "low";

dffeas \mem[5][57] (
	.clk(clk),
	.d(ShiftLeft157),
	.asdata(\mem[6][57]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][57]~q ),
	.prn(vcc));
defparam \mem[5][57] .is_wysiwyg = "true";
defparam \mem[5][57] .power_up = "low";

dffeas \mem[4][57] (
	.clk(clk),
	.d(ShiftLeft157),
	.asdata(\mem[5][57]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][57]~q ),
	.prn(vcc));
defparam \mem[4][57] .is_wysiwyg = "true";
defparam \mem[4][57] .power_up = "low";

dffeas \mem[3][57] (
	.clk(clk),
	.d(ShiftLeft157),
	.asdata(\mem[4][57]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][57]~q ),
	.prn(vcc));
defparam \mem[3][57] .is_wysiwyg = "true";
defparam \mem[3][57] .power_up = "low";

dffeas \mem[2][57] (
	.clk(clk),
	.d(ShiftLeft157),
	.asdata(\mem[3][57]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][57]~q ),
	.prn(vcc));
defparam \mem[2][57] .is_wysiwyg = "true";
defparam \mem[2][57] .power_up = "low";

dffeas \mem[1][57] (
	.clk(clk),
	.d(ShiftLeft157),
	.asdata(\mem[2][57]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][57]~q ),
	.prn(vcc));
defparam \mem[1][57] .is_wysiwyg = "true";
defparam \mem[1][57] .power_up = "low";

dffeas \mem[7][1] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][1]~q ),
	.prn(vcc));
defparam \mem[7][1] .is_wysiwyg = "true";
defparam \mem[7][1] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft11),
	.datac(!\mem[7][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h2727272727272727;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[6][1] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][1]~q ),
	.prn(vcc));
defparam \mem[6][1] .is_wysiwyg = "true";
defparam \mem[6][1] .power_up = "low";

dffeas \mem[5][1] (
	.clk(clk),
	.d(ShiftLeft11),
	.asdata(\mem[6][1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][1]~q ),
	.prn(vcc));
defparam \mem[5][1] .is_wysiwyg = "true";
defparam \mem[5][1] .power_up = "low";

dffeas \mem[4][1] (
	.clk(clk),
	.d(ShiftLeft11),
	.asdata(\mem[5][1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][1]~q ),
	.prn(vcc));
defparam \mem[4][1] .is_wysiwyg = "true";
defparam \mem[4][1] .power_up = "low";

dffeas \mem[3][1] (
	.clk(clk),
	.d(ShiftLeft11),
	.asdata(\mem[4][1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][1]~q ),
	.prn(vcc));
defparam \mem[3][1] .is_wysiwyg = "true";
defparam \mem[3][1] .power_up = "low";

dffeas \mem[2][1] (
	.clk(clk),
	.d(ShiftLeft11),
	.asdata(\mem[3][1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][1]~q ),
	.prn(vcc));
defparam \mem[2][1] .is_wysiwyg = "true";
defparam \mem[2][1] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(ShiftLeft11),
	.asdata(\mem[2][1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

dffeas \mem[7][33] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][33]~q ),
	.prn(vcc));
defparam \mem[7][33] .is_wysiwyg = "true";
defparam \mem[7][33] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft133),
	.datac(!\mem[7][33]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h2727272727272727;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[6][33] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][33]~q ),
	.prn(vcc));
defparam \mem[6][33] .is_wysiwyg = "true";
defparam \mem[6][33] .power_up = "low";

dffeas \mem[5][33] (
	.clk(clk),
	.d(ShiftLeft133),
	.asdata(\mem[6][33]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][33]~q ),
	.prn(vcc));
defparam \mem[5][33] .is_wysiwyg = "true";
defparam \mem[5][33] .power_up = "low";

dffeas \mem[4][33] (
	.clk(clk),
	.d(ShiftLeft133),
	.asdata(\mem[5][33]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][33]~q ),
	.prn(vcc));
defparam \mem[4][33] .is_wysiwyg = "true";
defparam \mem[4][33] .power_up = "low";

dffeas \mem[3][33] (
	.clk(clk),
	.d(ShiftLeft133),
	.asdata(\mem[4][33]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][33]~q ),
	.prn(vcc));
defparam \mem[3][33] .is_wysiwyg = "true";
defparam \mem[3][33] .power_up = "low";

dffeas \mem[2][33] (
	.clk(clk),
	.d(ShiftLeft133),
	.asdata(\mem[3][33]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][33]~q ),
	.prn(vcc));
defparam \mem[2][33] .is_wysiwyg = "true";
defparam \mem[2][33] .power_up = "low";

dffeas \mem[1][33] (
	.clk(clk),
	.d(ShiftLeft133),
	.asdata(\mem[2][33]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][33]~q ),
	.prn(vcc));
defparam \mem[1][33] .is_wysiwyg = "true";
defparam \mem[1][33] .power_up = "low";

dffeas \mem[7][10] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][10]~q ),
	.prn(vcc));
defparam \mem[7][10] .is_wysiwyg = "true";
defparam \mem[7][10] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft110),
	.datac(!\mem[7][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h2727272727272727;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[6][10] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][10]~q ),
	.prn(vcc));
defparam \mem[6][10] .is_wysiwyg = "true";
defparam \mem[6][10] .power_up = "low";

dffeas \mem[5][10] (
	.clk(clk),
	.d(ShiftLeft110),
	.asdata(\mem[6][10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][10]~q ),
	.prn(vcc));
defparam \mem[5][10] .is_wysiwyg = "true";
defparam \mem[5][10] .power_up = "low";

dffeas \mem[4][10] (
	.clk(clk),
	.d(ShiftLeft110),
	.asdata(\mem[5][10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][10]~q ),
	.prn(vcc));
defparam \mem[4][10] .is_wysiwyg = "true";
defparam \mem[4][10] .power_up = "low";

dffeas \mem[3][10] (
	.clk(clk),
	.d(ShiftLeft110),
	.asdata(\mem[4][10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][10]~q ),
	.prn(vcc));
defparam \mem[3][10] .is_wysiwyg = "true";
defparam \mem[3][10] .power_up = "low";

dffeas \mem[2][10] (
	.clk(clk),
	.d(ShiftLeft110),
	.asdata(\mem[3][10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][10]~q ),
	.prn(vcc));
defparam \mem[2][10] .is_wysiwyg = "true";
defparam \mem[2][10] .power_up = "low";

dffeas \mem[1][10] (
	.clk(clk),
	.d(ShiftLeft110),
	.asdata(\mem[2][10]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

dffeas \mem[7][42] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][42]~q ),
	.prn(vcc));
defparam \mem[7][42] .is_wysiwyg = "true";
defparam \mem[7][42] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft142),
	.datac(!\mem[7][42]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h2727272727272727;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[6][42] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][42]~q ),
	.prn(vcc));
defparam \mem[6][42] .is_wysiwyg = "true";
defparam \mem[6][42] .power_up = "low";

dffeas \mem[5][42] (
	.clk(clk),
	.d(ShiftLeft142),
	.asdata(\mem[6][42]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][42]~q ),
	.prn(vcc));
defparam \mem[5][42] .is_wysiwyg = "true";
defparam \mem[5][42] .power_up = "low";

dffeas \mem[4][42] (
	.clk(clk),
	.d(ShiftLeft142),
	.asdata(\mem[5][42]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][42]~q ),
	.prn(vcc));
defparam \mem[4][42] .is_wysiwyg = "true";
defparam \mem[4][42] .power_up = "low";

dffeas \mem[3][42] (
	.clk(clk),
	.d(ShiftLeft142),
	.asdata(\mem[4][42]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][42]~q ),
	.prn(vcc));
defparam \mem[3][42] .is_wysiwyg = "true";
defparam \mem[3][42] .power_up = "low";

dffeas \mem[2][42] (
	.clk(clk),
	.d(ShiftLeft142),
	.asdata(\mem[3][42]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][42]~q ),
	.prn(vcc));
defparam \mem[2][42] .is_wysiwyg = "true";
defparam \mem[2][42] .power_up = "low";

dffeas \mem[1][42] (
	.clk(clk),
	.d(ShiftLeft142),
	.asdata(\mem[2][42]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][42]~q ),
	.prn(vcc));
defparam \mem[1][42] .is_wysiwyg = "true";
defparam \mem[1][42] .power_up = "low";

dffeas \mem[7][18] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][18]~q ),
	.prn(vcc));
defparam \mem[7][18] .is_wysiwyg = "true";
defparam \mem[7][18] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft118),
	.datac(!\mem[7][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h2727272727272727;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[6][18] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][18]~q ),
	.prn(vcc));
defparam \mem[6][18] .is_wysiwyg = "true";
defparam \mem[6][18] .power_up = "low";

dffeas \mem[5][18] (
	.clk(clk),
	.d(ShiftLeft118),
	.asdata(\mem[6][18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][18]~q ),
	.prn(vcc));
defparam \mem[5][18] .is_wysiwyg = "true";
defparam \mem[5][18] .power_up = "low";

dffeas \mem[4][18] (
	.clk(clk),
	.d(ShiftLeft118),
	.asdata(\mem[5][18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][18]~q ),
	.prn(vcc));
defparam \mem[4][18] .is_wysiwyg = "true";
defparam \mem[4][18] .power_up = "low";

dffeas \mem[3][18] (
	.clk(clk),
	.d(ShiftLeft118),
	.asdata(\mem[4][18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][18]~q ),
	.prn(vcc));
defparam \mem[3][18] .is_wysiwyg = "true";
defparam \mem[3][18] .power_up = "low";

dffeas \mem[2][18] (
	.clk(clk),
	.d(ShiftLeft118),
	.asdata(\mem[3][18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][18]~q ),
	.prn(vcc));
defparam \mem[2][18] .is_wysiwyg = "true";
defparam \mem[2][18] .power_up = "low";

dffeas \mem[1][18] (
	.clk(clk),
	.d(ShiftLeft118),
	.asdata(\mem[2][18]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

dffeas \mem[7][50] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][50]~q ),
	.prn(vcc));
defparam \mem[7][50] .is_wysiwyg = "true";
defparam \mem[7][50] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft150),
	.datac(!\mem[7][50]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h2727272727272727;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[6][50] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][50]~q ),
	.prn(vcc));
defparam \mem[6][50] .is_wysiwyg = "true";
defparam \mem[6][50] .power_up = "low";

dffeas \mem[5][50] (
	.clk(clk),
	.d(ShiftLeft150),
	.asdata(\mem[6][50]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][50]~q ),
	.prn(vcc));
defparam \mem[5][50] .is_wysiwyg = "true";
defparam \mem[5][50] .power_up = "low";

dffeas \mem[4][50] (
	.clk(clk),
	.d(ShiftLeft150),
	.asdata(\mem[5][50]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][50]~q ),
	.prn(vcc));
defparam \mem[4][50] .is_wysiwyg = "true";
defparam \mem[4][50] .power_up = "low";

dffeas \mem[3][50] (
	.clk(clk),
	.d(ShiftLeft150),
	.asdata(\mem[4][50]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][50]~q ),
	.prn(vcc));
defparam \mem[3][50] .is_wysiwyg = "true";
defparam \mem[3][50] .power_up = "low";

dffeas \mem[2][50] (
	.clk(clk),
	.d(ShiftLeft150),
	.asdata(\mem[3][50]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][50]~q ),
	.prn(vcc));
defparam \mem[2][50] .is_wysiwyg = "true";
defparam \mem[2][50] .power_up = "low";

dffeas \mem[1][50] (
	.clk(clk),
	.d(ShiftLeft150),
	.asdata(\mem[2][50]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][50]~q ),
	.prn(vcc));
defparam \mem[1][50] .is_wysiwyg = "true";
defparam \mem[1][50] .power_up = "low";

dffeas \mem[7][26] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][26]~q ),
	.prn(vcc));
defparam \mem[7][26] .is_wysiwyg = "true";
defparam \mem[7][26] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft126),
	.datac(!\mem[7][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h2727272727272727;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[6][26] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][26]~q ),
	.prn(vcc));
defparam \mem[6][26] .is_wysiwyg = "true";
defparam \mem[6][26] .power_up = "low";

dffeas \mem[5][26] (
	.clk(clk),
	.d(ShiftLeft126),
	.asdata(\mem[6][26]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][26]~q ),
	.prn(vcc));
defparam \mem[5][26] .is_wysiwyg = "true";
defparam \mem[5][26] .power_up = "low";

dffeas \mem[4][26] (
	.clk(clk),
	.d(ShiftLeft126),
	.asdata(\mem[5][26]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][26]~q ),
	.prn(vcc));
defparam \mem[4][26] .is_wysiwyg = "true";
defparam \mem[4][26] .power_up = "low";

dffeas \mem[3][26] (
	.clk(clk),
	.d(ShiftLeft126),
	.asdata(\mem[4][26]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][26]~q ),
	.prn(vcc));
defparam \mem[3][26] .is_wysiwyg = "true";
defparam \mem[3][26] .power_up = "low";

dffeas \mem[2][26] (
	.clk(clk),
	.d(ShiftLeft126),
	.asdata(\mem[3][26]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][26]~q ),
	.prn(vcc));
defparam \mem[2][26] .is_wysiwyg = "true";
defparam \mem[2][26] .power_up = "low";

dffeas \mem[1][26] (
	.clk(clk),
	.d(ShiftLeft126),
	.asdata(\mem[2][26]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

dffeas \mem[7][58] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][58]~q ),
	.prn(vcc));
defparam \mem[7][58] .is_wysiwyg = "true";
defparam \mem[7][58] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft158),
	.datac(!\mem[7][58]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h2727272727272727;
defparam \mem~31 .shared_arith = "off";

dffeas \mem[6][58] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][58]~q ),
	.prn(vcc));
defparam \mem[6][58] .is_wysiwyg = "true";
defparam \mem[6][58] .power_up = "low";

dffeas \mem[5][58] (
	.clk(clk),
	.d(ShiftLeft158),
	.asdata(\mem[6][58]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][58]~q ),
	.prn(vcc));
defparam \mem[5][58] .is_wysiwyg = "true";
defparam \mem[5][58] .power_up = "low";

dffeas \mem[4][58] (
	.clk(clk),
	.d(ShiftLeft158),
	.asdata(\mem[5][58]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][58]~q ),
	.prn(vcc));
defparam \mem[4][58] .is_wysiwyg = "true";
defparam \mem[4][58] .power_up = "low";

dffeas \mem[3][58] (
	.clk(clk),
	.d(ShiftLeft158),
	.asdata(\mem[4][58]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][58]~q ),
	.prn(vcc));
defparam \mem[3][58] .is_wysiwyg = "true";
defparam \mem[3][58] .power_up = "low";

dffeas \mem[2][58] (
	.clk(clk),
	.d(ShiftLeft158),
	.asdata(\mem[3][58]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][58]~q ),
	.prn(vcc));
defparam \mem[2][58] .is_wysiwyg = "true";
defparam \mem[2][58] .power_up = "low";

dffeas \mem[1][58] (
	.clk(clk),
	.d(ShiftLeft158),
	.asdata(\mem[2][58]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][58]~q ),
	.prn(vcc));
defparam \mem[1][58] .is_wysiwyg = "true";
defparam \mem[1][58] .power_up = "low";

dffeas \mem[7][2] (
	.clk(clk),
	.d(\mem~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][2]~q ),
	.prn(vcc));
defparam \mem[7][2] .is_wysiwyg = "true";
defparam \mem[7][2] .power_up = "low";

cyclonev_lcell_comb \mem~32 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft12),
	.datac(!\mem[7][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~32 .extended_lut = "off";
defparam \mem~32 .lut_mask = 64'h2727272727272727;
defparam \mem~32 .shared_arith = "off";

dffeas \mem[6][2] (
	.clk(clk),
	.d(\mem~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][2]~q ),
	.prn(vcc));
defparam \mem[6][2] .is_wysiwyg = "true";
defparam \mem[6][2] .power_up = "low";

dffeas \mem[5][2] (
	.clk(clk),
	.d(ShiftLeft12),
	.asdata(\mem[6][2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][2]~q ),
	.prn(vcc));
defparam \mem[5][2] .is_wysiwyg = "true";
defparam \mem[5][2] .power_up = "low";

dffeas \mem[4][2] (
	.clk(clk),
	.d(ShiftLeft12),
	.asdata(\mem[5][2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][2]~q ),
	.prn(vcc));
defparam \mem[4][2] .is_wysiwyg = "true";
defparam \mem[4][2] .power_up = "low";

dffeas \mem[3][2] (
	.clk(clk),
	.d(ShiftLeft12),
	.asdata(\mem[4][2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][2]~q ),
	.prn(vcc));
defparam \mem[3][2] .is_wysiwyg = "true";
defparam \mem[3][2] .power_up = "low";

dffeas \mem[2][2] (
	.clk(clk),
	.d(ShiftLeft12),
	.asdata(\mem[3][2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][2]~q ),
	.prn(vcc));
defparam \mem[2][2] .is_wysiwyg = "true";
defparam \mem[2][2] .power_up = "low";

dffeas \mem[1][2] (
	.clk(clk),
	.d(ShiftLeft12),
	.asdata(\mem[2][2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

dffeas \mem[7][34] (
	.clk(clk),
	.d(\mem~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][34]~q ),
	.prn(vcc));
defparam \mem[7][34] .is_wysiwyg = "true";
defparam \mem[7][34] .power_up = "low";

cyclonev_lcell_comb \mem~33 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft134),
	.datac(!\mem[7][34]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~33 .extended_lut = "off";
defparam \mem~33 .lut_mask = 64'h2727272727272727;
defparam \mem~33 .shared_arith = "off";

dffeas \mem[6][34] (
	.clk(clk),
	.d(\mem~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][34]~q ),
	.prn(vcc));
defparam \mem[6][34] .is_wysiwyg = "true";
defparam \mem[6][34] .power_up = "low";

dffeas \mem[5][34] (
	.clk(clk),
	.d(ShiftLeft134),
	.asdata(\mem[6][34]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][34]~q ),
	.prn(vcc));
defparam \mem[5][34] .is_wysiwyg = "true";
defparam \mem[5][34] .power_up = "low";

dffeas \mem[4][34] (
	.clk(clk),
	.d(ShiftLeft134),
	.asdata(\mem[5][34]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][34]~q ),
	.prn(vcc));
defparam \mem[4][34] .is_wysiwyg = "true";
defparam \mem[4][34] .power_up = "low";

dffeas \mem[3][34] (
	.clk(clk),
	.d(ShiftLeft134),
	.asdata(\mem[4][34]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][34]~q ),
	.prn(vcc));
defparam \mem[3][34] .is_wysiwyg = "true";
defparam \mem[3][34] .power_up = "low";

dffeas \mem[2][34] (
	.clk(clk),
	.d(ShiftLeft134),
	.asdata(\mem[3][34]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][34]~q ),
	.prn(vcc));
defparam \mem[2][34] .is_wysiwyg = "true";
defparam \mem[2][34] .power_up = "low";

dffeas \mem[1][34] (
	.clk(clk),
	.d(ShiftLeft134),
	.asdata(\mem[2][34]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][34]~q ),
	.prn(vcc));
defparam \mem[1][34] .is_wysiwyg = "true";
defparam \mem[1][34] .power_up = "low";

dffeas \mem[7][11] (
	.clk(clk),
	.d(\mem~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][11]~q ),
	.prn(vcc));
defparam \mem[7][11] .is_wysiwyg = "true";
defparam \mem[7][11] .power_up = "low";

cyclonev_lcell_comb \mem~34 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft111),
	.datac(!\mem[7][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~34 .extended_lut = "off";
defparam \mem~34 .lut_mask = 64'h2727272727272727;
defparam \mem~34 .shared_arith = "off";

dffeas \mem[6][11] (
	.clk(clk),
	.d(\mem~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][11]~q ),
	.prn(vcc));
defparam \mem[6][11] .is_wysiwyg = "true";
defparam \mem[6][11] .power_up = "low";

dffeas \mem[5][11] (
	.clk(clk),
	.d(ShiftLeft111),
	.asdata(\mem[6][11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][11]~q ),
	.prn(vcc));
defparam \mem[5][11] .is_wysiwyg = "true";
defparam \mem[5][11] .power_up = "low";

dffeas \mem[4][11] (
	.clk(clk),
	.d(ShiftLeft111),
	.asdata(\mem[5][11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][11]~q ),
	.prn(vcc));
defparam \mem[4][11] .is_wysiwyg = "true";
defparam \mem[4][11] .power_up = "low";

dffeas \mem[3][11] (
	.clk(clk),
	.d(ShiftLeft111),
	.asdata(\mem[4][11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][11]~q ),
	.prn(vcc));
defparam \mem[3][11] .is_wysiwyg = "true";
defparam \mem[3][11] .power_up = "low";

dffeas \mem[2][11] (
	.clk(clk),
	.d(ShiftLeft111),
	.asdata(\mem[3][11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][11]~q ),
	.prn(vcc));
defparam \mem[2][11] .is_wysiwyg = "true";
defparam \mem[2][11] .power_up = "low";

dffeas \mem[1][11] (
	.clk(clk),
	.d(ShiftLeft111),
	.asdata(\mem[2][11]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

dffeas \mem[7][43] (
	.clk(clk),
	.d(\mem~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][43]~q ),
	.prn(vcc));
defparam \mem[7][43] .is_wysiwyg = "true";
defparam \mem[7][43] .power_up = "low";

cyclonev_lcell_comb \mem~35 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft143),
	.datac(!\mem[7][43]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~35 .extended_lut = "off";
defparam \mem~35 .lut_mask = 64'h2727272727272727;
defparam \mem~35 .shared_arith = "off";

dffeas \mem[6][43] (
	.clk(clk),
	.d(\mem~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][43]~q ),
	.prn(vcc));
defparam \mem[6][43] .is_wysiwyg = "true";
defparam \mem[6][43] .power_up = "low";

dffeas \mem[5][43] (
	.clk(clk),
	.d(ShiftLeft143),
	.asdata(\mem[6][43]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][43]~q ),
	.prn(vcc));
defparam \mem[5][43] .is_wysiwyg = "true";
defparam \mem[5][43] .power_up = "low";

dffeas \mem[4][43] (
	.clk(clk),
	.d(ShiftLeft143),
	.asdata(\mem[5][43]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][43]~q ),
	.prn(vcc));
defparam \mem[4][43] .is_wysiwyg = "true";
defparam \mem[4][43] .power_up = "low";

dffeas \mem[3][43] (
	.clk(clk),
	.d(ShiftLeft143),
	.asdata(\mem[4][43]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][43]~q ),
	.prn(vcc));
defparam \mem[3][43] .is_wysiwyg = "true";
defparam \mem[3][43] .power_up = "low";

dffeas \mem[2][43] (
	.clk(clk),
	.d(ShiftLeft143),
	.asdata(\mem[3][43]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][43]~q ),
	.prn(vcc));
defparam \mem[2][43] .is_wysiwyg = "true";
defparam \mem[2][43] .power_up = "low";

dffeas \mem[1][43] (
	.clk(clk),
	.d(ShiftLeft143),
	.asdata(\mem[2][43]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][43]~q ),
	.prn(vcc));
defparam \mem[1][43] .is_wysiwyg = "true";
defparam \mem[1][43] .power_up = "low";

dffeas \mem[7][19] (
	.clk(clk),
	.d(\mem~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][19]~q ),
	.prn(vcc));
defparam \mem[7][19] .is_wysiwyg = "true";
defparam \mem[7][19] .power_up = "low";

cyclonev_lcell_comb \mem~36 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft119),
	.datac(!\mem[7][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~36 .extended_lut = "off";
defparam \mem~36 .lut_mask = 64'h2727272727272727;
defparam \mem~36 .shared_arith = "off";

dffeas \mem[6][19] (
	.clk(clk),
	.d(\mem~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][19]~q ),
	.prn(vcc));
defparam \mem[6][19] .is_wysiwyg = "true";
defparam \mem[6][19] .power_up = "low";

dffeas \mem[5][19] (
	.clk(clk),
	.d(ShiftLeft119),
	.asdata(\mem[6][19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][19]~q ),
	.prn(vcc));
defparam \mem[5][19] .is_wysiwyg = "true";
defparam \mem[5][19] .power_up = "low";

dffeas \mem[4][19] (
	.clk(clk),
	.d(ShiftLeft119),
	.asdata(\mem[5][19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][19]~q ),
	.prn(vcc));
defparam \mem[4][19] .is_wysiwyg = "true";
defparam \mem[4][19] .power_up = "low";

dffeas \mem[3][19] (
	.clk(clk),
	.d(ShiftLeft119),
	.asdata(\mem[4][19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][19]~q ),
	.prn(vcc));
defparam \mem[3][19] .is_wysiwyg = "true";
defparam \mem[3][19] .power_up = "low";

dffeas \mem[2][19] (
	.clk(clk),
	.d(ShiftLeft119),
	.asdata(\mem[3][19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][19]~q ),
	.prn(vcc));
defparam \mem[2][19] .is_wysiwyg = "true";
defparam \mem[2][19] .power_up = "low";

dffeas \mem[1][19] (
	.clk(clk),
	.d(ShiftLeft119),
	.asdata(\mem[2][19]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

dffeas \mem[7][51] (
	.clk(clk),
	.d(\mem~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][51]~q ),
	.prn(vcc));
defparam \mem[7][51] .is_wysiwyg = "true";
defparam \mem[7][51] .power_up = "low";

cyclonev_lcell_comb \mem~37 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft151),
	.datac(!\mem[7][51]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~37 .extended_lut = "off";
defparam \mem~37 .lut_mask = 64'h2727272727272727;
defparam \mem~37 .shared_arith = "off";

dffeas \mem[6][51] (
	.clk(clk),
	.d(\mem~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][51]~q ),
	.prn(vcc));
defparam \mem[6][51] .is_wysiwyg = "true";
defparam \mem[6][51] .power_up = "low";

dffeas \mem[5][51] (
	.clk(clk),
	.d(ShiftLeft151),
	.asdata(\mem[6][51]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][51]~q ),
	.prn(vcc));
defparam \mem[5][51] .is_wysiwyg = "true";
defparam \mem[5][51] .power_up = "low";

dffeas \mem[4][51] (
	.clk(clk),
	.d(ShiftLeft151),
	.asdata(\mem[5][51]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][51]~q ),
	.prn(vcc));
defparam \mem[4][51] .is_wysiwyg = "true";
defparam \mem[4][51] .power_up = "low";

dffeas \mem[3][51] (
	.clk(clk),
	.d(ShiftLeft151),
	.asdata(\mem[4][51]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][51]~q ),
	.prn(vcc));
defparam \mem[3][51] .is_wysiwyg = "true";
defparam \mem[3][51] .power_up = "low";

dffeas \mem[2][51] (
	.clk(clk),
	.d(ShiftLeft151),
	.asdata(\mem[3][51]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][51]~q ),
	.prn(vcc));
defparam \mem[2][51] .is_wysiwyg = "true";
defparam \mem[2][51] .power_up = "low";

dffeas \mem[1][51] (
	.clk(clk),
	.d(ShiftLeft151),
	.asdata(\mem[2][51]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][51]~q ),
	.prn(vcc));
defparam \mem[1][51] .is_wysiwyg = "true";
defparam \mem[1][51] .power_up = "low";

dffeas \mem[7][27] (
	.clk(clk),
	.d(\mem~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][27]~q ),
	.prn(vcc));
defparam \mem[7][27] .is_wysiwyg = "true";
defparam \mem[7][27] .power_up = "low";

cyclonev_lcell_comb \mem~38 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft127),
	.datac(!\mem[7][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~38 .extended_lut = "off";
defparam \mem~38 .lut_mask = 64'h2727272727272727;
defparam \mem~38 .shared_arith = "off";

dffeas \mem[6][27] (
	.clk(clk),
	.d(\mem~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][27]~q ),
	.prn(vcc));
defparam \mem[6][27] .is_wysiwyg = "true";
defparam \mem[6][27] .power_up = "low";

dffeas \mem[5][27] (
	.clk(clk),
	.d(ShiftLeft127),
	.asdata(\mem[6][27]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][27]~q ),
	.prn(vcc));
defparam \mem[5][27] .is_wysiwyg = "true";
defparam \mem[5][27] .power_up = "low";

dffeas \mem[4][27] (
	.clk(clk),
	.d(ShiftLeft127),
	.asdata(\mem[5][27]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][27]~q ),
	.prn(vcc));
defparam \mem[4][27] .is_wysiwyg = "true";
defparam \mem[4][27] .power_up = "low";

dffeas \mem[3][27] (
	.clk(clk),
	.d(ShiftLeft127),
	.asdata(\mem[4][27]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][27]~q ),
	.prn(vcc));
defparam \mem[3][27] .is_wysiwyg = "true";
defparam \mem[3][27] .power_up = "low";

dffeas \mem[2][27] (
	.clk(clk),
	.d(ShiftLeft127),
	.asdata(\mem[3][27]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][27]~q ),
	.prn(vcc));
defparam \mem[2][27] .is_wysiwyg = "true";
defparam \mem[2][27] .power_up = "low";

dffeas \mem[1][27] (
	.clk(clk),
	.d(ShiftLeft127),
	.asdata(\mem[2][27]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

dffeas \mem[7][59] (
	.clk(clk),
	.d(\mem~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][59]~q ),
	.prn(vcc));
defparam \mem[7][59] .is_wysiwyg = "true";
defparam \mem[7][59] .power_up = "low";

cyclonev_lcell_comb \mem~39 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft159),
	.datac(!\mem[7][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~39 .extended_lut = "off";
defparam \mem~39 .lut_mask = 64'h2727272727272727;
defparam \mem~39 .shared_arith = "off";

dffeas \mem[6][59] (
	.clk(clk),
	.d(\mem~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][59]~q ),
	.prn(vcc));
defparam \mem[6][59] .is_wysiwyg = "true";
defparam \mem[6][59] .power_up = "low";

dffeas \mem[5][59] (
	.clk(clk),
	.d(ShiftLeft159),
	.asdata(\mem[6][59]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][59]~q ),
	.prn(vcc));
defparam \mem[5][59] .is_wysiwyg = "true";
defparam \mem[5][59] .power_up = "low";

dffeas \mem[4][59] (
	.clk(clk),
	.d(ShiftLeft159),
	.asdata(\mem[5][59]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][59]~q ),
	.prn(vcc));
defparam \mem[4][59] .is_wysiwyg = "true";
defparam \mem[4][59] .power_up = "low";

dffeas \mem[3][59] (
	.clk(clk),
	.d(ShiftLeft159),
	.asdata(\mem[4][59]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][59]~q ),
	.prn(vcc));
defparam \mem[3][59] .is_wysiwyg = "true";
defparam \mem[3][59] .power_up = "low";

dffeas \mem[2][59] (
	.clk(clk),
	.d(ShiftLeft159),
	.asdata(\mem[3][59]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][59]~q ),
	.prn(vcc));
defparam \mem[2][59] .is_wysiwyg = "true";
defparam \mem[2][59] .power_up = "low";

dffeas \mem[1][59] (
	.clk(clk),
	.d(ShiftLeft159),
	.asdata(\mem[2][59]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

dffeas \mem[7][3] (
	.clk(clk),
	.d(\mem~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][3]~q ),
	.prn(vcc));
defparam \mem[7][3] .is_wysiwyg = "true";
defparam \mem[7][3] .power_up = "low";

cyclonev_lcell_comb \mem~40 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft13),
	.datac(!\mem[7][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~40 .extended_lut = "off";
defparam \mem~40 .lut_mask = 64'h2727272727272727;
defparam \mem~40 .shared_arith = "off";

dffeas \mem[6][3] (
	.clk(clk),
	.d(\mem~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][3]~q ),
	.prn(vcc));
defparam \mem[6][3] .is_wysiwyg = "true";
defparam \mem[6][3] .power_up = "low";

dffeas \mem[5][3] (
	.clk(clk),
	.d(ShiftLeft13),
	.asdata(\mem[6][3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][3]~q ),
	.prn(vcc));
defparam \mem[5][3] .is_wysiwyg = "true";
defparam \mem[5][3] .power_up = "low";

dffeas \mem[4][3] (
	.clk(clk),
	.d(ShiftLeft13),
	.asdata(\mem[5][3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][3]~q ),
	.prn(vcc));
defparam \mem[4][3] .is_wysiwyg = "true";
defparam \mem[4][3] .power_up = "low";

dffeas \mem[3][3] (
	.clk(clk),
	.d(ShiftLeft13),
	.asdata(\mem[4][3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][3]~q ),
	.prn(vcc));
defparam \mem[3][3] .is_wysiwyg = "true";
defparam \mem[3][3] .power_up = "low";

dffeas \mem[2][3] (
	.clk(clk),
	.d(ShiftLeft13),
	.asdata(\mem[3][3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][3]~q ),
	.prn(vcc));
defparam \mem[2][3] .is_wysiwyg = "true";
defparam \mem[2][3] .power_up = "low";

dffeas \mem[1][3] (
	.clk(clk),
	.d(ShiftLeft13),
	.asdata(\mem[2][3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

dffeas \mem[7][35] (
	.clk(clk),
	.d(\mem~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][35]~q ),
	.prn(vcc));
defparam \mem[7][35] .is_wysiwyg = "true";
defparam \mem[7][35] .power_up = "low";

cyclonev_lcell_comb \mem~41 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft135),
	.datac(!\mem[7][35]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~41 .extended_lut = "off";
defparam \mem~41 .lut_mask = 64'h2727272727272727;
defparam \mem~41 .shared_arith = "off";

dffeas \mem[6][35] (
	.clk(clk),
	.d(\mem~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][35]~q ),
	.prn(vcc));
defparam \mem[6][35] .is_wysiwyg = "true";
defparam \mem[6][35] .power_up = "low";

dffeas \mem[5][35] (
	.clk(clk),
	.d(ShiftLeft135),
	.asdata(\mem[6][35]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][35]~q ),
	.prn(vcc));
defparam \mem[5][35] .is_wysiwyg = "true";
defparam \mem[5][35] .power_up = "low";

dffeas \mem[4][35] (
	.clk(clk),
	.d(ShiftLeft135),
	.asdata(\mem[5][35]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][35]~q ),
	.prn(vcc));
defparam \mem[4][35] .is_wysiwyg = "true";
defparam \mem[4][35] .power_up = "low";

dffeas \mem[3][35] (
	.clk(clk),
	.d(ShiftLeft135),
	.asdata(\mem[4][35]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][35]~q ),
	.prn(vcc));
defparam \mem[3][35] .is_wysiwyg = "true";
defparam \mem[3][35] .power_up = "low";

dffeas \mem[2][35] (
	.clk(clk),
	.d(ShiftLeft135),
	.asdata(\mem[3][35]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][35]~q ),
	.prn(vcc));
defparam \mem[2][35] .is_wysiwyg = "true";
defparam \mem[2][35] .power_up = "low";

dffeas \mem[1][35] (
	.clk(clk),
	.d(ShiftLeft135),
	.asdata(\mem[2][35]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][35]~q ),
	.prn(vcc));
defparam \mem[1][35] .is_wysiwyg = "true";
defparam \mem[1][35] .power_up = "low";

dffeas \mem[7][12] (
	.clk(clk),
	.d(\mem~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][12]~q ),
	.prn(vcc));
defparam \mem[7][12] .is_wysiwyg = "true";
defparam \mem[7][12] .power_up = "low";

cyclonev_lcell_comb \mem~42 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft112),
	.datac(!\mem[7][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~42 .extended_lut = "off";
defparam \mem~42 .lut_mask = 64'h2727272727272727;
defparam \mem~42 .shared_arith = "off";

dffeas \mem[6][12] (
	.clk(clk),
	.d(\mem~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][12]~q ),
	.prn(vcc));
defparam \mem[6][12] .is_wysiwyg = "true";
defparam \mem[6][12] .power_up = "low";

dffeas \mem[5][12] (
	.clk(clk),
	.d(ShiftLeft112),
	.asdata(\mem[6][12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][12]~q ),
	.prn(vcc));
defparam \mem[5][12] .is_wysiwyg = "true";
defparam \mem[5][12] .power_up = "low";

dffeas \mem[4][12] (
	.clk(clk),
	.d(ShiftLeft112),
	.asdata(\mem[5][12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][12]~q ),
	.prn(vcc));
defparam \mem[4][12] .is_wysiwyg = "true";
defparam \mem[4][12] .power_up = "low";

dffeas \mem[3][12] (
	.clk(clk),
	.d(ShiftLeft112),
	.asdata(\mem[4][12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][12]~q ),
	.prn(vcc));
defparam \mem[3][12] .is_wysiwyg = "true";
defparam \mem[3][12] .power_up = "low";

dffeas \mem[2][12] (
	.clk(clk),
	.d(ShiftLeft112),
	.asdata(\mem[3][12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][12]~q ),
	.prn(vcc));
defparam \mem[2][12] .is_wysiwyg = "true";
defparam \mem[2][12] .power_up = "low";

dffeas \mem[1][12] (
	.clk(clk),
	.d(ShiftLeft112),
	.asdata(\mem[2][12]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

dffeas \mem[7][44] (
	.clk(clk),
	.d(\mem~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][44]~q ),
	.prn(vcc));
defparam \mem[7][44] .is_wysiwyg = "true";
defparam \mem[7][44] .power_up = "low";

cyclonev_lcell_comb \mem~43 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft144),
	.datac(!\mem[7][44]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~43 .extended_lut = "off";
defparam \mem~43 .lut_mask = 64'h2727272727272727;
defparam \mem~43 .shared_arith = "off";

dffeas \mem[6][44] (
	.clk(clk),
	.d(\mem~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][44]~q ),
	.prn(vcc));
defparam \mem[6][44] .is_wysiwyg = "true";
defparam \mem[6][44] .power_up = "low";

dffeas \mem[5][44] (
	.clk(clk),
	.d(ShiftLeft144),
	.asdata(\mem[6][44]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][44]~q ),
	.prn(vcc));
defparam \mem[5][44] .is_wysiwyg = "true";
defparam \mem[5][44] .power_up = "low";

dffeas \mem[4][44] (
	.clk(clk),
	.d(ShiftLeft144),
	.asdata(\mem[5][44]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][44]~q ),
	.prn(vcc));
defparam \mem[4][44] .is_wysiwyg = "true";
defparam \mem[4][44] .power_up = "low";

dffeas \mem[3][44] (
	.clk(clk),
	.d(ShiftLeft144),
	.asdata(\mem[4][44]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][44]~q ),
	.prn(vcc));
defparam \mem[3][44] .is_wysiwyg = "true";
defparam \mem[3][44] .power_up = "low";

dffeas \mem[2][44] (
	.clk(clk),
	.d(ShiftLeft144),
	.asdata(\mem[3][44]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][44]~q ),
	.prn(vcc));
defparam \mem[2][44] .is_wysiwyg = "true";
defparam \mem[2][44] .power_up = "low";

dffeas \mem[1][44] (
	.clk(clk),
	.d(ShiftLeft144),
	.asdata(\mem[2][44]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][44]~q ),
	.prn(vcc));
defparam \mem[1][44] .is_wysiwyg = "true";
defparam \mem[1][44] .power_up = "low";

dffeas \mem[7][20] (
	.clk(clk),
	.d(\mem~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][20]~q ),
	.prn(vcc));
defparam \mem[7][20] .is_wysiwyg = "true";
defparam \mem[7][20] .power_up = "low";

cyclonev_lcell_comb \mem~44 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft120),
	.datac(!\mem[7][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~44 .extended_lut = "off";
defparam \mem~44 .lut_mask = 64'h2727272727272727;
defparam \mem~44 .shared_arith = "off";

dffeas \mem[6][20] (
	.clk(clk),
	.d(\mem~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][20]~q ),
	.prn(vcc));
defparam \mem[6][20] .is_wysiwyg = "true";
defparam \mem[6][20] .power_up = "low";

dffeas \mem[5][20] (
	.clk(clk),
	.d(ShiftLeft120),
	.asdata(\mem[6][20]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][20]~q ),
	.prn(vcc));
defparam \mem[5][20] .is_wysiwyg = "true";
defparam \mem[5][20] .power_up = "low";

dffeas \mem[4][20] (
	.clk(clk),
	.d(ShiftLeft120),
	.asdata(\mem[5][20]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][20]~q ),
	.prn(vcc));
defparam \mem[4][20] .is_wysiwyg = "true";
defparam \mem[4][20] .power_up = "low";

dffeas \mem[3][20] (
	.clk(clk),
	.d(ShiftLeft120),
	.asdata(\mem[4][20]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][20]~q ),
	.prn(vcc));
defparam \mem[3][20] .is_wysiwyg = "true";
defparam \mem[3][20] .power_up = "low";

dffeas \mem[2][20] (
	.clk(clk),
	.d(ShiftLeft120),
	.asdata(\mem[3][20]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][20]~q ),
	.prn(vcc));
defparam \mem[2][20] .is_wysiwyg = "true";
defparam \mem[2][20] .power_up = "low";

dffeas \mem[1][20] (
	.clk(clk),
	.d(ShiftLeft120),
	.asdata(\mem[2][20]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

dffeas \mem[7][52] (
	.clk(clk),
	.d(\mem~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][52]~q ),
	.prn(vcc));
defparam \mem[7][52] .is_wysiwyg = "true";
defparam \mem[7][52] .power_up = "low";

cyclonev_lcell_comb \mem~45 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft152),
	.datac(!\mem[7][52]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~45 .extended_lut = "off";
defparam \mem~45 .lut_mask = 64'h2727272727272727;
defparam \mem~45 .shared_arith = "off";

dffeas \mem[6][52] (
	.clk(clk),
	.d(\mem~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][52]~q ),
	.prn(vcc));
defparam \mem[6][52] .is_wysiwyg = "true";
defparam \mem[6][52] .power_up = "low";

dffeas \mem[5][52] (
	.clk(clk),
	.d(ShiftLeft152),
	.asdata(\mem[6][52]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][52]~q ),
	.prn(vcc));
defparam \mem[5][52] .is_wysiwyg = "true";
defparam \mem[5][52] .power_up = "low";

dffeas \mem[4][52] (
	.clk(clk),
	.d(ShiftLeft152),
	.asdata(\mem[5][52]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][52]~q ),
	.prn(vcc));
defparam \mem[4][52] .is_wysiwyg = "true";
defparam \mem[4][52] .power_up = "low";

dffeas \mem[3][52] (
	.clk(clk),
	.d(ShiftLeft152),
	.asdata(\mem[4][52]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][52]~q ),
	.prn(vcc));
defparam \mem[3][52] .is_wysiwyg = "true";
defparam \mem[3][52] .power_up = "low";

dffeas \mem[2][52] (
	.clk(clk),
	.d(ShiftLeft152),
	.asdata(\mem[3][52]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][52]~q ),
	.prn(vcc));
defparam \mem[2][52] .is_wysiwyg = "true";
defparam \mem[2][52] .power_up = "low";

dffeas \mem[1][52] (
	.clk(clk),
	.d(ShiftLeft152),
	.asdata(\mem[2][52]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][52]~q ),
	.prn(vcc));
defparam \mem[1][52] .is_wysiwyg = "true";
defparam \mem[1][52] .power_up = "low";

dffeas \mem[7][28] (
	.clk(clk),
	.d(\mem~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][28]~q ),
	.prn(vcc));
defparam \mem[7][28] .is_wysiwyg = "true";
defparam \mem[7][28] .power_up = "low";

cyclonev_lcell_comb \mem~46 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft128),
	.datac(!\mem[7][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~46 .extended_lut = "off";
defparam \mem~46 .lut_mask = 64'h2727272727272727;
defparam \mem~46 .shared_arith = "off";

dffeas \mem[6][28] (
	.clk(clk),
	.d(\mem~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][28]~q ),
	.prn(vcc));
defparam \mem[6][28] .is_wysiwyg = "true";
defparam \mem[6][28] .power_up = "low";

dffeas \mem[5][28] (
	.clk(clk),
	.d(ShiftLeft128),
	.asdata(\mem[6][28]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][28]~q ),
	.prn(vcc));
defparam \mem[5][28] .is_wysiwyg = "true";
defparam \mem[5][28] .power_up = "low";

dffeas \mem[4][28] (
	.clk(clk),
	.d(ShiftLeft128),
	.asdata(\mem[5][28]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][28]~q ),
	.prn(vcc));
defparam \mem[4][28] .is_wysiwyg = "true";
defparam \mem[4][28] .power_up = "low";

dffeas \mem[3][28] (
	.clk(clk),
	.d(ShiftLeft128),
	.asdata(\mem[4][28]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][28]~q ),
	.prn(vcc));
defparam \mem[3][28] .is_wysiwyg = "true";
defparam \mem[3][28] .power_up = "low";

dffeas \mem[2][28] (
	.clk(clk),
	.d(ShiftLeft128),
	.asdata(\mem[3][28]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][28]~q ),
	.prn(vcc));
defparam \mem[2][28] .is_wysiwyg = "true";
defparam \mem[2][28] .power_up = "low";

dffeas \mem[1][28] (
	.clk(clk),
	.d(ShiftLeft128),
	.asdata(\mem[2][28]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

dffeas \mem[7][60] (
	.clk(clk),
	.d(\mem~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][60]~q ),
	.prn(vcc));
defparam \mem[7][60] .is_wysiwyg = "true";
defparam \mem[7][60] .power_up = "low";

cyclonev_lcell_comb \mem~47 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft160),
	.datac(!\mem[7][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~47 .extended_lut = "off";
defparam \mem~47 .lut_mask = 64'h2727272727272727;
defparam \mem~47 .shared_arith = "off";

dffeas \mem[6][60] (
	.clk(clk),
	.d(\mem~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][60]~q ),
	.prn(vcc));
defparam \mem[6][60] .is_wysiwyg = "true";
defparam \mem[6][60] .power_up = "low";

dffeas \mem[5][60] (
	.clk(clk),
	.d(ShiftLeft160),
	.asdata(\mem[6][60]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][60]~q ),
	.prn(vcc));
defparam \mem[5][60] .is_wysiwyg = "true";
defparam \mem[5][60] .power_up = "low";

dffeas \mem[4][60] (
	.clk(clk),
	.d(ShiftLeft160),
	.asdata(\mem[5][60]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][60]~q ),
	.prn(vcc));
defparam \mem[4][60] .is_wysiwyg = "true";
defparam \mem[4][60] .power_up = "low";

dffeas \mem[3][60] (
	.clk(clk),
	.d(ShiftLeft160),
	.asdata(\mem[4][60]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][60]~q ),
	.prn(vcc));
defparam \mem[3][60] .is_wysiwyg = "true";
defparam \mem[3][60] .power_up = "low";

dffeas \mem[2][60] (
	.clk(clk),
	.d(ShiftLeft160),
	.asdata(\mem[3][60]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][60]~q ),
	.prn(vcc));
defparam \mem[2][60] .is_wysiwyg = "true";
defparam \mem[2][60] .power_up = "low";

dffeas \mem[1][60] (
	.clk(clk),
	.d(ShiftLeft160),
	.asdata(\mem[2][60]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

dffeas \mem[7][4] (
	.clk(clk),
	.d(\mem~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][4]~q ),
	.prn(vcc));
defparam \mem[7][4] .is_wysiwyg = "true";
defparam \mem[7][4] .power_up = "low";

cyclonev_lcell_comb \mem~48 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft14),
	.datac(!\mem[7][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~48 .extended_lut = "off";
defparam \mem~48 .lut_mask = 64'h2727272727272727;
defparam \mem~48 .shared_arith = "off";

dffeas \mem[6][4] (
	.clk(clk),
	.d(\mem~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][4]~q ),
	.prn(vcc));
defparam \mem[6][4] .is_wysiwyg = "true";
defparam \mem[6][4] .power_up = "low";

dffeas \mem[5][4] (
	.clk(clk),
	.d(ShiftLeft14),
	.asdata(\mem[6][4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][4]~q ),
	.prn(vcc));
defparam \mem[5][4] .is_wysiwyg = "true";
defparam \mem[5][4] .power_up = "low";

dffeas \mem[4][4] (
	.clk(clk),
	.d(ShiftLeft14),
	.asdata(\mem[5][4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][4]~q ),
	.prn(vcc));
defparam \mem[4][4] .is_wysiwyg = "true";
defparam \mem[4][4] .power_up = "low";

dffeas \mem[3][4] (
	.clk(clk),
	.d(ShiftLeft14),
	.asdata(\mem[4][4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][4]~q ),
	.prn(vcc));
defparam \mem[3][4] .is_wysiwyg = "true";
defparam \mem[3][4] .power_up = "low";

dffeas \mem[2][4] (
	.clk(clk),
	.d(ShiftLeft14),
	.asdata(\mem[3][4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][4]~q ),
	.prn(vcc));
defparam \mem[2][4] .is_wysiwyg = "true";
defparam \mem[2][4] .power_up = "low";

dffeas \mem[1][4] (
	.clk(clk),
	.d(ShiftLeft14),
	.asdata(\mem[2][4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

dffeas \mem[7][36] (
	.clk(clk),
	.d(\mem~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][36]~q ),
	.prn(vcc));
defparam \mem[7][36] .is_wysiwyg = "true";
defparam \mem[7][36] .power_up = "low";

cyclonev_lcell_comb \mem~49 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft136),
	.datac(!\mem[7][36]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~49 .extended_lut = "off";
defparam \mem~49 .lut_mask = 64'h2727272727272727;
defparam \mem~49 .shared_arith = "off";

dffeas \mem[6][36] (
	.clk(clk),
	.d(\mem~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][36]~q ),
	.prn(vcc));
defparam \mem[6][36] .is_wysiwyg = "true";
defparam \mem[6][36] .power_up = "low";

dffeas \mem[5][36] (
	.clk(clk),
	.d(ShiftLeft136),
	.asdata(\mem[6][36]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][36]~q ),
	.prn(vcc));
defparam \mem[5][36] .is_wysiwyg = "true";
defparam \mem[5][36] .power_up = "low";

dffeas \mem[4][36] (
	.clk(clk),
	.d(ShiftLeft136),
	.asdata(\mem[5][36]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][36]~q ),
	.prn(vcc));
defparam \mem[4][36] .is_wysiwyg = "true";
defparam \mem[4][36] .power_up = "low";

dffeas \mem[3][36] (
	.clk(clk),
	.d(ShiftLeft136),
	.asdata(\mem[4][36]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][36]~q ),
	.prn(vcc));
defparam \mem[3][36] .is_wysiwyg = "true";
defparam \mem[3][36] .power_up = "low";

dffeas \mem[2][36] (
	.clk(clk),
	.d(ShiftLeft136),
	.asdata(\mem[3][36]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][36]~q ),
	.prn(vcc));
defparam \mem[2][36] .is_wysiwyg = "true";
defparam \mem[2][36] .power_up = "low";

dffeas \mem[1][36] (
	.clk(clk),
	.d(ShiftLeft136),
	.asdata(\mem[2][36]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][36]~q ),
	.prn(vcc));
defparam \mem[1][36] .is_wysiwyg = "true";
defparam \mem[1][36] .power_up = "low";

dffeas \mem[7][13] (
	.clk(clk),
	.d(\mem~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][13]~q ),
	.prn(vcc));
defparam \mem[7][13] .is_wysiwyg = "true";
defparam \mem[7][13] .power_up = "low";

cyclonev_lcell_comb \mem~50 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft113),
	.datac(!\mem[7][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~50 .extended_lut = "off";
defparam \mem~50 .lut_mask = 64'h2727272727272727;
defparam \mem~50 .shared_arith = "off";

dffeas \mem[6][13] (
	.clk(clk),
	.d(\mem~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][13]~q ),
	.prn(vcc));
defparam \mem[6][13] .is_wysiwyg = "true";
defparam \mem[6][13] .power_up = "low";

dffeas \mem[5][13] (
	.clk(clk),
	.d(ShiftLeft113),
	.asdata(\mem[6][13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][13]~q ),
	.prn(vcc));
defparam \mem[5][13] .is_wysiwyg = "true";
defparam \mem[5][13] .power_up = "low";

dffeas \mem[4][13] (
	.clk(clk),
	.d(ShiftLeft113),
	.asdata(\mem[5][13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][13]~q ),
	.prn(vcc));
defparam \mem[4][13] .is_wysiwyg = "true";
defparam \mem[4][13] .power_up = "low";

dffeas \mem[3][13] (
	.clk(clk),
	.d(ShiftLeft113),
	.asdata(\mem[4][13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][13]~q ),
	.prn(vcc));
defparam \mem[3][13] .is_wysiwyg = "true";
defparam \mem[3][13] .power_up = "low";

dffeas \mem[2][13] (
	.clk(clk),
	.d(ShiftLeft113),
	.asdata(\mem[3][13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][13]~q ),
	.prn(vcc));
defparam \mem[2][13] .is_wysiwyg = "true";
defparam \mem[2][13] .power_up = "low";

dffeas \mem[1][13] (
	.clk(clk),
	.d(ShiftLeft113),
	.asdata(\mem[2][13]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

dffeas \mem[7][45] (
	.clk(clk),
	.d(\mem~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][45]~q ),
	.prn(vcc));
defparam \mem[7][45] .is_wysiwyg = "true";
defparam \mem[7][45] .power_up = "low";

cyclonev_lcell_comb \mem~51 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft145),
	.datac(!\mem[7][45]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~51 .extended_lut = "off";
defparam \mem~51 .lut_mask = 64'h2727272727272727;
defparam \mem~51 .shared_arith = "off";

dffeas \mem[6][45] (
	.clk(clk),
	.d(\mem~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][45]~q ),
	.prn(vcc));
defparam \mem[6][45] .is_wysiwyg = "true";
defparam \mem[6][45] .power_up = "low";

dffeas \mem[5][45] (
	.clk(clk),
	.d(ShiftLeft145),
	.asdata(\mem[6][45]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][45]~q ),
	.prn(vcc));
defparam \mem[5][45] .is_wysiwyg = "true";
defparam \mem[5][45] .power_up = "low";

dffeas \mem[4][45] (
	.clk(clk),
	.d(ShiftLeft145),
	.asdata(\mem[5][45]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][45]~q ),
	.prn(vcc));
defparam \mem[4][45] .is_wysiwyg = "true";
defparam \mem[4][45] .power_up = "low";

dffeas \mem[3][45] (
	.clk(clk),
	.d(ShiftLeft145),
	.asdata(\mem[4][45]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][45]~q ),
	.prn(vcc));
defparam \mem[3][45] .is_wysiwyg = "true";
defparam \mem[3][45] .power_up = "low";

dffeas \mem[2][45] (
	.clk(clk),
	.d(ShiftLeft145),
	.asdata(\mem[3][45]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][45]~q ),
	.prn(vcc));
defparam \mem[2][45] .is_wysiwyg = "true";
defparam \mem[2][45] .power_up = "low";

dffeas \mem[1][45] (
	.clk(clk),
	.d(ShiftLeft145),
	.asdata(\mem[2][45]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][45]~q ),
	.prn(vcc));
defparam \mem[1][45] .is_wysiwyg = "true";
defparam \mem[1][45] .power_up = "low";

dffeas \mem[7][21] (
	.clk(clk),
	.d(\mem~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][21]~q ),
	.prn(vcc));
defparam \mem[7][21] .is_wysiwyg = "true";
defparam \mem[7][21] .power_up = "low";

cyclonev_lcell_comb \mem~52 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft121),
	.datac(!\mem[7][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~52 .extended_lut = "off";
defparam \mem~52 .lut_mask = 64'h2727272727272727;
defparam \mem~52 .shared_arith = "off";

dffeas \mem[6][21] (
	.clk(clk),
	.d(\mem~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][21]~q ),
	.prn(vcc));
defparam \mem[6][21] .is_wysiwyg = "true";
defparam \mem[6][21] .power_up = "low";

dffeas \mem[5][21] (
	.clk(clk),
	.d(ShiftLeft121),
	.asdata(\mem[6][21]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][21]~q ),
	.prn(vcc));
defparam \mem[5][21] .is_wysiwyg = "true";
defparam \mem[5][21] .power_up = "low";

dffeas \mem[4][21] (
	.clk(clk),
	.d(ShiftLeft121),
	.asdata(\mem[5][21]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][21]~q ),
	.prn(vcc));
defparam \mem[4][21] .is_wysiwyg = "true";
defparam \mem[4][21] .power_up = "low";

dffeas \mem[3][21] (
	.clk(clk),
	.d(ShiftLeft121),
	.asdata(\mem[4][21]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][21]~q ),
	.prn(vcc));
defparam \mem[3][21] .is_wysiwyg = "true";
defparam \mem[3][21] .power_up = "low";

dffeas \mem[2][21] (
	.clk(clk),
	.d(ShiftLeft121),
	.asdata(\mem[3][21]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][21]~q ),
	.prn(vcc));
defparam \mem[2][21] .is_wysiwyg = "true";
defparam \mem[2][21] .power_up = "low";

dffeas \mem[1][21] (
	.clk(clk),
	.d(ShiftLeft121),
	.asdata(\mem[2][21]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

dffeas \mem[7][53] (
	.clk(clk),
	.d(\mem~53_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][53]~q ),
	.prn(vcc));
defparam \mem[7][53] .is_wysiwyg = "true";
defparam \mem[7][53] .power_up = "low";

cyclonev_lcell_comb \mem~53 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft153),
	.datac(!\mem[7][53]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~53 .extended_lut = "off";
defparam \mem~53 .lut_mask = 64'h2727272727272727;
defparam \mem~53 .shared_arith = "off";

dffeas \mem[6][53] (
	.clk(clk),
	.d(\mem~53_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][53]~q ),
	.prn(vcc));
defparam \mem[6][53] .is_wysiwyg = "true";
defparam \mem[6][53] .power_up = "low";

dffeas \mem[5][53] (
	.clk(clk),
	.d(ShiftLeft153),
	.asdata(\mem[6][53]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][53]~q ),
	.prn(vcc));
defparam \mem[5][53] .is_wysiwyg = "true";
defparam \mem[5][53] .power_up = "low";

dffeas \mem[4][53] (
	.clk(clk),
	.d(ShiftLeft153),
	.asdata(\mem[5][53]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][53]~q ),
	.prn(vcc));
defparam \mem[4][53] .is_wysiwyg = "true";
defparam \mem[4][53] .power_up = "low";

dffeas \mem[3][53] (
	.clk(clk),
	.d(ShiftLeft153),
	.asdata(\mem[4][53]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][53]~q ),
	.prn(vcc));
defparam \mem[3][53] .is_wysiwyg = "true";
defparam \mem[3][53] .power_up = "low";

dffeas \mem[2][53] (
	.clk(clk),
	.d(ShiftLeft153),
	.asdata(\mem[3][53]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][53]~q ),
	.prn(vcc));
defparam \mem[2][53] .is_wysiwyg = "true";
defparam \mem[2][53] .power_up = "low";

dffeas \mem[1][53] (
	.clk(clk),
	.d(ShiftLeft153),
	.asdata(\mem[2][53]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][53]~q ),
	.prn(vcc));
defparam \mem[1][53] .is_wysiwyg = "true";
defparam \mem[1][53] .power_up = "low";

dffeas \mem[7][29] (
	.clk(clk),
	.d(\mem~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][29]~q ),
	.prn(vcc));
defparam \mem[7][29] .is_wysiwyg = "true";
defparam \mem[7][29] .power_up = "low";

cyclonev_lcell_comb \mem~54 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft129),
	.datac(!\mem[7][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~54 .extended_lut = "off";
defparam \mem~54 .lut_mask = 64'h2727272727272727;
defparam \mem~54 .shared_arith = "off";

dffeas \mem[6][29] (
	.clk(clk),
	.d(\mem~54_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][29]~q ),
	.prn(vcc));
defparam \mem[6][29] .is_wysiwyg = "true";
defparam \mem[6][29] .power_up = "low";

dffeas \mem[5][29] (
	.clk(clk),
	.d(ShiftLeft129),
	.asdata(\mem[6][29]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][29]~q ),
	.prn(vcc));
defparam \mem[5][29] .is_wysiwyg = "true";
defparam \mem[5][29] .power_up = "low";

dffeas \mem[4][29] (
	.clk(clk),
	.d(ShiftLeft129),
	.asdata(\mem[5][29]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][29]~q ),
	.prn(vcc));
defparam \mem[4][29] .is_wysiwyg = "true";
defparam \mem[4][29] .power_up = "low";

dffeas \mem[3][29] (
	.clk(clk),
	.d(ShiftLeft129),
	.asdata(\mem[4][29]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][29]~q ),
	.prn(vcc));
defparam \mem[3][29] .is_wysiwyg = "true";
defparam \mem[3][29] .power_up = "low";

dffeas \mem[2][29] (
	.clk(clk),
	.d(ShiftLeft129),
	.asdata(\mem[3][29]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][29]~q ),
	.prn(vcc));
defparam \mem[2][29] .is_wysiwyg = "true";
defparam \mem[2][29] .power_up = "low";

dffeas \mem[1][29] (
	.clk(clk),
	.d(ShiftLeft129),
	.asdata(\mem[2][29]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

dffeas \mem[7][61] (
	.clk(clk),
	.d(\mem~55_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][61]~q ),
	.prn(vcc));
defparam \mem[7][61] .is_wysiwyg = "true";
defparam \mem[7][61] .power_up = "low";

cyclonev_lcell_comb \mem~55 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft161),
	.datac(!\mem[7][61]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~55 .extended_lut = "off";
defparam \mem~55 .lut_mask = 64'h2727272727272727;
defparam \mem~55 .shared_arith = "off";

dffeas \mem[6][61] (
	.clk(clk),
	.d(\mem~55_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][61]~q ),
	.prn(vcc));
defparam \mem[6][61] .is_wysiwyg = "true";
defparam \mem[6][61] .power_up = "low";

dffeas \mem[5][61] (
	.clk(clk),
	.d(ShiftLeft161),
	.asdata(\mem[6][61]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][61]~q ),
	.prn(vcc));
defparam \mem[5][61] .is_wysiwyg = "true";
defparam \mem[5][61] .power_up = "low";

dffeas \mem[4][61] (
	.clk(clk),
	.d(ShiftLeft161),
	.asdata(\mem[5][61]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][61]~q ),
	.prn(vcc));
defparam \mem[4][61] .is_wysiwyg = "true";
defparam \mem[4][61] .power_up = "low";

dffeas \mem[3][61] (
	.clk(clk),
	.d(ShiftLeft161),
	.asdata(\mem[4][61]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][61]~q ),
	.prn(vcc));
defparam \mem[3][61] .is_wysiwyg = "true";
defparam \mem[3][61] .power_up = "low";

dffeas \mem[2][61] (
	.clk(clk),
	.d(ShiftLeft161),
	.asdata(\mem[3][61]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][61]~q ),
	.prn(vcc));
defparam \mem[2][61] .is_wysiwyg = "true";
defparam \mem[2][61] .power_up = "low";

dffeas \mem[1][61] (
	.clk(clk),
	.d(ShiftLeft161),
	.asdata(\mem[2][61]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][61]~q ),
	.prn(vcc));
defparam \mem[1][61] .is_wysiwyg = "true";
defparam \mem[1][61] .power_up = "low";

dffeas \mem[7][5] (
	.clk(clk),
	.d(\mem~56_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][5]~q ),
	.prn(vcc));
defparam \mem[7][5] .is_wysiwyg = "true";
defparam \mem[7][5] .power_up = "low";

cyclonev_lcell_comb \mem~56 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft15),
	.datac(!\mem[7][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~56 .extended_lut = "off";
defparam \mem~56 .lut_mask = 64'h2727272727272727;
defparam \mem~56 .shared_arith = "off";

dffeas \mem[6][5] (
	.clk(clk),
	.d(\mem~56_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][5]~q ),
	.prn(vcc));
defparam \mem[6][5] .is_wysiwyg = "true";
defparam \mem[6][5] .power_up = "low";

dffeas \mem[5][5] (
	.clk(clk),
	.d(ShiftLeft15),
	.asdata(\mem[6][5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][5]~q ),
	.prn(vcc));
defparam \mem[5][5] .is_wysiwyg = "true";
defparam \mem[5][5] .power_up = "low";

dffeas \mem[4][5] (
	.clk(clk),
	.d(ShiftLeft15),
	.asdata(\mem[5][5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][5]~q ),
	.prn(vcc));
defparam \mem[4][5] .is_wysiwyg = "true";
defparam \mem[4][5] .power_up = "low";

dffeas \mem[3][5] (
	.clk(clk),
	.d(ShiftLeft15),
	.asdata(\mem[4][5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][5]~q ),
	.prn(vcc));
defparam \mem[3][5] .is_wysiwyg = "true";
defparam \mem[3][5] .power_up = "low";

dffeas \mem[2][5] (
	.clk(clk),
	.d(ShiftLeft15),
	.asdata(\mem[3][5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][5]~q ),
	.prn(vcc));
defparam \mem[2][5] .is_wysiwyg = "true";
defparam \mem[2][5] .power_up = "low";

dffeas \mem[1][5] (
	.clk(clk),
	.d(ShiftLeft15),
	.asdata(\mem[2][5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

dffeas \mem[7][37] (
	.clk(clk),
	.d(\mem~57_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][37]~q ),
	.prn(vcc));
defparam \mem[7][37] .is_wysiwyg = "true";
defparam \mem[7][37] .power_up = "low";

cyclonev_lcell_comb \mem~57 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft137),
	.datac(!\mem[7][37]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~57 .extended_lut = "off";
defparam \mem~57 .lut_mask = 64'h2727272727272727;
defparam \mem~57 .shared_arith = "off";

dffeas \mem[6][37] (
	.clk(clk),
	.d(\mem~57_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][37]~q ),
	.prn(vcc));
defparam \mem[6][37] .is_wysiwyg = "true";
defparam \mem[6][37] .power_up = "low";

dffeas \mem[5][37] (
	.clk(clk),
	.d(ShiftLeft137),
	.asdata(\mem[6][37]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][37]~q ),
	.prn(vcc));
defparam \mem[5][37] .is_wysiwyg = "true";
defparam \mem[5][37] .power_up = "low";

dffeas \mem[4][37] (
	.clk(clk),
	.d(ShiftLeft137),
	.asdata(\mem[5][37]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][37]~q ),
	.prn(vcc));
defparam \mem[4][37] .is_wysiwyg = "true";
defparam \mem[4][37] .power_up = "low";

dffeas \mem[3][37] (
	.clk(clk),
	.d(ShiftLeft137),
	.asdata(\mem[4][37]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][37]~q ),
	.prn(vcc));
defparam \mem[3][37] .is_wysiwyg = "true";
defparam \mem[3][37] .power_up = "low";

dffeas \mem[2][37] (
	.clk(clk),
	.d(ShiftLeft137),
	.asdata(\mem[3][37]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][37]~q ),
	.prn(vcc));
defparam \mem[2][37] .is_wysiwyg = "true";
defparam \mem[2][37] .power_up = "low";

dffeas \mem[1][37] (
	.clk(clk),
	.d(ShiftLeft137),
	.asdata(\mem[2][37]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][37]~q ),
	.prn(vcc));
defparam \mem[1][37] .is_wysiwyg = "true";
defparam \mem[1][37] .power_up = "low";

dffeas \mem[7][14] (
	.clk(clk),
	.d(\mem~58_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][14]~q ),
	.prn(vcc));
defparam \mem[7][14] .is_wysiwyg = "true";
defparam \mem[7][14] .power_up = "low";

cyclonev_lcell_comb \mem~58 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft114),
	.datac(!\mem[7][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~58 .extended_lut = "off";
defparam \mem~58 .lut_mask = 64'h2727272727272727;
defparam \mem~58 .shared_arith = "off";

dffeas \mem[6][14] (
	.clk(clk),
	.d(\mem~58_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][14]~q ),
	.prn(vcc));
defparam \mem[6][14] .is_wysiwyg = "true";
defparam \mem[6][14] .power_up = "low";

dffeas \mem[5][14] (
	.clk(clk),
	.d(ShiftLeft114),
	.asdata(\mem[6][14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][14]~q ),
	.prn(vcc));
defparam \mem[5][14] .is_wysiwyg = "true";
defparam \mem[5][14] .power_up = "low";

dffeas \mem[4][14] (
	.clk(clk),
	.d(ShiftLeft114),
	.asdata(\mem[5][14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][14]~q ),
	.prn(vcc));
defparam \mem[4][14] .is_wysiwyg = "true";
defparam \mem[4][14] .power_up = "low";

dffeas \mem[3][14] (
	.clk(clk),
	.d(ShiftLeft114),
	.asdata(\mem[4][14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][14]~q ),
	.prn(vcc));
defparam \mem[3][14] .is_wysiwyg = "true";
defparam \mem[3][14] .power_up = "low";

dffeas \mem[2][14] (
	.clk(clk),
	.d(ShiftLeft114),
	.asdata(\mem[3][14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][14]~q ),
	.prn(vcc));
defparam \mem[2][14] .is_wysiwyg = "true";
defparam \mem[2][14] .power_up = "low";

dffeas \mem[1][14] (
	.clk(clk),
	.d(ShiftLeft114),
	.asdata(\mem[2][14]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

dffeas \mem[7][46] (
	.clk(clk),
	.d(\mem~59_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][46]~q ),
	.prn(vcc));
defparam \mem[7][46] .is_wysiwyg = "true";
defparam \mem[7][46] .power_up = "low";

cyclonev_lcell_comb \mem~59 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft146),
	.datac(!\mem[7][46]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~59 .extended_lut = "off";
defparam \mem~59 .lut_mask = 64'h2727272727272727;
defparam \mem~59 .shared_arith = "off";

dffeas \mem[6][46] (
	.clk(clk),
	.d(\mem~59_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][46]~q ),
	.prn(vcc));
defparam \mem[6][46] .is_wysiwyg = "true";
defparam \mem[6][46] .power_up = "low";

dffeas \mem[5][46] (
	.clk(clk),
	.d(ShiftLeft146),
	.asdata(\mem[6][46]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][46]~q ),
	.prn(vcc));
defparam \mem[5][46] .is_wysiwyg = "true";
defparam \mem[5][46] .power_up = "low";

dffeas \mem[4][46] (
	.clk(clk),
	.d(ShiftLeft146),
	.asdata(\mem[5][46]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][46]~q ),
	.prn(vcc));
defparam \mem[4][46] .is_wysiwyg = "true";
defparam \mem[4][46] .power_up = "low";

dffeas \mem[3][46] (
	.clk(clk),
	.d(ShiftLeft146),
	.asdata(\mem[4][46]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][46]~q ),
	.prn(vcc));
defparam \mem[3][46] .is_wysiwyg = "true";
defparam \mem[3][46] .power_up = "low";

dffeas \mem[2][46] (
	.clk(clk),
	.d(ShiftLeft146),
	.asdata(\mem[3][46]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][46]~q ),
	.prn(vcc));
defparam \mem[2][46] .is_wysiwyg = "true";
defparam \mem[2][46] .power_up = "low";

dffeas \mem[1][46] (
	.clk(clk),
	.d(ShiftLeft146),
	.asdata(\mem[2][46]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][46]~q ),
	.prn(vcc));
defparam \mem[1][46] .is_wysiwyg = "true";
defparam \mem[1][46] .power_up = "low";

dffeas \mem[7][22] (
	.clk(clk),
	.d(\mem~60_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][22]~q ),
	.prn(vcc));
defparam \mem[7][22] .is_wysiwyg = "true";
defparam \mem[7][22] .power_up = "low";

cyclonev_lcell_comb \mem~60 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft122),
	.datac(!\mem[7][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~60 .extended_lut = "off";
defparam \mem~60 .lut_mask = 64'h2727272727272727;
defparam \mem~60 .shared_arith = "off";

dffeas \mem[6][22] (
	.clk(clk),
	.d(\mem~60_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][22]~q ),
	.prn(vcc));
defparam \mem[6][22] .is_wysiwyg = "true";
defparam \mem[6][22] .power_up = "low";

dffeas \mem[5][22] (
	.clk(clk),
	.d(ShiftLeft122),
	.asdata(\mem[6][22]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][22]~q ),
	.prn(vcc));
defparam \mem[5][22] .is_wysiwyg = "true";
defparam \mem[5][22] .power_up = "low";

dffeas \mem[4][22] (
	.clk(clk),
	.d(ShiftLeft122),
	.asdata(\mem[5][22]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][22]~q ),
	.prn(vcc));
defparam \mem[4][22] .is_wysiwyg = "true";
defparam \mem[4][22] .power_up = "low";

dffeas \mem[3][22] (
	.clk(clk),
	.d(ShiftLeft122),
	.asdata(\mem[4][22]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][22]~q ),
	.prn(vcc));
defparam \mem[3][22] .is_wysiwyg = "true";
defparam \mem[3][22] .power_up = "low";

dffeas \mem[2][22] (
	.clk(clk),
	.d(ShiftLeft122),
	.asdata(\mem[3][22]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][22]~q ),
	.prn(vcc));
defparam \mem[2][22] .is_wysiwyg = "true";
defparam \mem[2][22] .power_up = "low";

dffeas \mem[1][22] (
	.clk(clk),
	.d(ShiftLeft122),
	.asdata(\mem[2][22]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

dffeas \mem[7][54] (
	.clk(clk),
	.d(\mem~61_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][54]~q ),
	.prn(vcc));
defparam \mem[7][54] .is_wysiwyg = "true";
defparam \mem[7][54] .power_up = "low";

cyclonev_lcell_comb \mem~61 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft154),
	.datac(!\mem[7][54]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~61 .extended_lut = "off";
defparam \mem~61 .lut_mask = 64'h2727272727272727;
defparam \mem~61 .shared_arith = "off";

dffeas \mem[6][54] (
	.clk(clk),
	.d(\mem~61_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][54]~q ),
	.prn(vcc));
defparam \mem[6][54] .is_wysiwyg = "true";
defparam \mem[6][54] .power_up = "low";

dffeas \mem[5][54] (
	.clk(clk),
	.d(ShiftLeft154),
	.asdata(\mem[6][54]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][54]~q ),
	.prn(vcc));
defparam \mem[5][54] .is_wysiwyg = "true";
defparam \mem[5][54] .power_up = "low";

dffeas \mem[4][54] (
	.clk(clk),
	.d(ShiftLeft154),
	.asdata(\mem[5][54]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][54]~q ),
	.prn(vcc));
defparam \mem[4][54] .is_wysiwyg = "true";
defparam \mem[4][54] .power_up = "low";

dffeas \mem[3][54] (
	.clk(clk),
	.d(ShiftLeft154),
	.asdata(\mem[4][54]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][54]~q ),
	.prn(vcc));
defparam \mem[3][54] .is_wysiwyg = "true";
defparam \mem[3][54] .power_up = "low";

dffeas \mem[2][54] (
	.clk(clk),
	.d(ShiftLeft154),
	.asdata(\mem[3][54]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][54]~q ),
	.prn(vcc));
defparam \mem[2][54] .is_wysiwyg = "true";
defparam \mem[2][54] .power_up = "low";

dffeas \mem[1][54] (
	.clk(clk),
	.d(ShiftLeft154),
	.asdata(\mem[2][54]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][54]~q ),
	.prn(vcc));
defparam \mem[1][54] .is_wysiwyg = "true";
defparam \mem[1][54] .power_up = "low";

dffeas \mem[7][30] (
	.clk(clk),
	.d(\mem~62_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][30]~q ),
	.prn(vcc));
defparam \mem[7][30] .is_wysiwyg = "true";
defparam \mem[7][30] .power_up = "low";

cyclonev_lcell_comb \mem~62 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft130),
	.datac(!\mem[7][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~62 .extended_lut = "off";
defparam \mem~62 .lut_mask = 64'h2727272727272727;
defparam \mem~62 .shared_arith = "off";

dffeas \mem[6][30] (
	.clk(clk),
	.d(\mem~62_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][30]~q ),
	.prn(vcc));
defparam \mem[6][30] .is_wysiwyg = "true";
defparam \mem[6][30] .power_up = "low";

dffeas \mem[5][30] (
	.clk(clk),
	.d(ShiftLeft130),
	.asdata(\mem[6][30]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][30]~q ),
	.prn(vcc));
defparam \mem[5][30] .is_wysiwyg = "true";
defparam \mem[5][30] .power_up = "low";

dffeas \mem[4][30] (
	.clk(clk),
	.d(ShiftLeft130),
	.asdata(\mem[5][30]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][30]~q ),
	.prn(vcc));
defparam \mem[4][30] .is_wysiwyg = "true";
defparam \mem[4][30] .power_up = "low";

dffeas \mem[3][30] (
	.clk(clk),
	.d(ShiftLeft130),
	.asdata(\mem[4][30]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][30]~q ),
	.prn(vcc));
defparam \mem[3][30] .is_wysiwyg = "true";
defparam \mem[3][30] .power_up = "low";

dffeas \mem[2][30] (
	.clk(clk),
	.d(ShiftLeft130),
	.asdata(\mem[3][30]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][30]~q ),
	.prn(vcc));
defparam \mem[2][30] .is_wysiwyg = "true";
defparam \mem[2][30] .power_up = "low";

dffeas \mem[1][30] (
	.clk(clk),
	.d(ShiftLeft130),
	.asdata(\mem[2][30]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

dffeas \mem[7][62] (
	.clk(clk),
	.d(\mem~63_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][62]~q ),
	.prn(vcc));
defparam \mem[7][62] .is_wysiwyg = "true";
defparam \mem[7][62] .power_up = "low";

cyclonev_lcell_comb \mem~63 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft162),
	.datac(!\mem[7][62]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~63 .extended_lut = "off";
defparam \mem~63 .lut_mask = 64'h2727272727272727;
defparam \mem~63 .shared_arith = "off";

dffeas \mem[6][62] (
	.clk(clk),
	.d(\mem~63_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][62]~q ),
	.prn(vcc));
defparam \mem[6][62] .is_wysiwyg = "true";
defparam \mem[6][62] .power_up = "low";

dffeas \mem[5][62] (
	.clk(clk),
	.d(ShiftLeft162),
	.asdata(\mem[6][62]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][62]~q ),
	.prn(vcc));
defparam \mem[5][62] .is_wysiwyg = "true";
defparam \mem[5][62] .power_up = "low";

dffeas \mem[4][62] (
	.clk(clk),
	.d(ShiftLeft162),
	.asdata(\mem[5][62]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][62]~q ),
	.prn(vcc));
defparam \mem[4][62] .is_wysiwyg = "true";
defparam \mem[4][62] .power_up = "low";

dffeas \mem[3][62] (
	.clk(clk),
	.d(ShiftLeft162),
	.asdata(\mem[4][62]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][62]~q ),
	.prn(vcc));
defparam \mem[3][62] .is_wysiwyg = "true";
defparam \mem[3][62] .power_up = "low";

dffeas \mem[2][62] (
	.clk(clk),
	.d(ShiftLeft162),
	.asdata(\mem[3][62]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][62]~q ),
	.prn(vcc));
defparam \mem[2][62] .is_wysiwyg = "true";
defparam \mem[2][62] .power_up = "low";

dffeas \mem[1][62] (
	.clk(clk),
	.d(ShiftLeft162),
	.asdata(\mem[2][62]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][62]~q ),
	.prn(vcc));
defparam \mem[1][62] .is_wysiwyg = "true";
defparam \mem[1][62] .power_up = "low";

dffeas \mem[7][6] (
	.clk(clk),
	.d(\mem~64_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][6]~q ),
	.prn(vcc));
defparam \mem[7][6] .is_wysiwyg = "true";
defparam \mem[7][6] .power_up = "low";

cyclonev_lcell_comb \mem~64 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft16),
	.datac(!\mem[7][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~64 .extended_lut = "off";
defparam \mem~64 .lut_mask = 64'h2727272727272727;
defparam \mem~64 .shared_arith = "off";

dffeas \mem[6][6] (
	.clk(clk),
	.d(\mem~64_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][6]~q ),
	.prn(vcc));
defparam \mem[6][6] .is_wysiwyg = "true";
defparam \mem[6][6] .power_up = "low";

dffeas \mem[5][6] (
	.clk(clk),
	.d(ShiftLeft16),
	.asdata(\mem[6][6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][6]~q ),
	.prn(vcc));
defparam \mem[5][6] .is_wysiwyg = "true";
defparam \mem[5][6] .power_up = "low";

dffeas \mem[4][6] (
	.clk(clk),
	.d(ShiftLeft16),
	.asdata(\mem[5][6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][6]~q ),
	.prn(vcc));
defparam \mem[4][6] .is_wysiwyg = "true";
defparam \mem[4][6] .power_up = "low";

dffeas \mem[3][6] (
	.clk(clk),
	.d(ShiftLeft16),
	.asdata(\mem[4][6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][6]~q ),
	.prn(vcc));
defparam \mem[3][6] .is_wysiwyg = "true";
defparam \mem[3][6] .power_up = "low";

dffeas \mem[2][6] (
	.clk(clk),
	.d(ShiftLeft16),
	.asdata(\mem[3][6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][6]~q ),
	.prn(vcc));
defparam \mem[2][6] .is_wysiwyg = "true";
defparam \mem[2][6] .power_up = "low";

dffeas \mem[1][6] (
	.clk(clk),
	.d(ShiftLeft16),
	.asdata(\mem[2][6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

dffeas \mem[7][38] (
	.clk(clk),
	.d(\mem~65_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][38]~q ),
	.prn(vcc));
defparam \mem[7][38] .is_wysiwyg = "true";
defparam \mem[7][38] .power_up = "low";

cyclonev_lcell_comb \mem~65 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft138),
	.datac(!\mem[7][38]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~65 .extended_lut = "off";
defparam \mem~65 .lut_mask = 64'h2727272727272727;
defparam \mem~65 .shared_arith = "off";

dffeas \mem[6][38] (
	.clk(clk),
	.d(\mem~65_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][38]~q ),
	.prn(vcc));
defparam \mem[6][38] .is_wysiwyg = "true";
defparam \mem[6][38] .power_up = "low";

dffeas \mem[5][38] (
	.clk(clk),
	.d(ShiftLeft138),
	.asdata(\mem[6][38]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][38]~q ),
	.prn(vcc));
defparam \mem[5][38] .is_wysiwyg = "true";
defparam \mem[5][38] .power_up = "low";

dffeas \mem[4][38] (
	.clk(clk),
	.d(ShiftLeft138),
	.asdata(\mem[5][38]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][38]~q ),
	.prn(vcc));
defparam \mem[4][38] .is_wysiwyg = "true";
defparam \mem[4][38] .power_up = "low";

dffeas \mem[3][38] (
	.clk(clk),
	.d(ShiftLeft138),
	.asdata(\mem[4][38]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][38]~q ),
	.prn(vcc));
defparam \mem[3][38] .is_wysiwyg = "true";
defparam \mem[3][38] .power_up = "low";

dffeas \mem[2][38] (
	.clk(clk),
	.d(ShiftLeft138),
	.asdata(\mem[3][38]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][38]~q ),
	.prn(vcc));
defparam \mem[2][38] .is_wysiwyg = "true";
defparam \mem[2][38] .power_up = "low";

dffeas \mem[1][38] (
	.clk(clk),
	.d(ShiftLeft138),
	.asdata(\mem[2][38]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][38]~q ),
	.prn(vcc));
defparam \mem[1][38] .is_wysiwyg = "true";
defparam \mem[1][38] .power_up = "low";

dffeas \mem[7][15] (
	.clk(clk),
	.d(\mem~66_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][15]~q ),
	.prn(vcc));
defparam \mem[7][15] .is_wysiwyg = "true";
defparam \mem[7][15] .power_up = "low";

cyclonev_lcell_comb \mem~66 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft115),
	.datac(!\mem[7][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~66 .extended_lut = "off";
defparam \mem~66 .lut_mask = 64'h2727272727272727;
defparam \mem~66 .shared_arith = "off";

dffeas \mem[6][15] (
	.clk(clk),
	.d(\mem~66_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][15]~q ),
	.prn(vcc));
defparam \mem[6][15] .is_wysiwyg = "true";
defparam \mem[6][15] .power_up = "low";

dffeas \mem[5][15] (
	.clk(clk),
	.d(ShiftLeft115),
	.asdata(\mem[6][15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][15]~q ),
	.prn(vcc));
defparam \mem[5][15] .is_wysiwyg = "true";
defparam \mem[5][15] .power_up = "low";

dffeas \mem[4][15] (
	.clk(clk),
	.d(ShiftLeft115),
	.asdata(\mem[5][15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][15]~q ),
	.prn(vcc));
defparam \mem[4][15] .is_wysiwyg = "true";
defparam \mem[4][15] .power_up = "low";

dffeas \mem[3][15] (
	.clk(clk),
	.d(ShiftLeft115),
	.asdata(\mem[4][15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][15]~q ),
	.prn(vcc));
defparam \mem[3][15] .is_wysiwyg = "true";
defparam \mem[3][15] .power_up = "low";

dffeas \mem[2][15] (
	.clk(clk),
	.d(ShiftLeft115),
	.asdata(\mem[3][15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][15]~q ),
	.prn(vcc));
defparam \mem[2][15] .is_wysiwyg = "true";
defparam \mem[2][15] .power_up = "low";

dffeas \mem[1][15] (
	.clk(clk),
	.d(ShiftLeft115),
	.asdata(\mem[2][15]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

dffeas \mem[7][47] (
	.clk(clk),
	.d(\mem~67_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][47]~q ),
	.prn(vcc));
defparam \mem[7][47] .is_wysiwyg = "true";
defparam \mem[7][47] .power_up = "low";

cyclonev_lcell_comb \mem~67 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft147),
	.datac(!\mem[7][47]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~67 .extended_lut = "off";
defparam \mem~67 .lut_mask = 64'h2727272727272727;
defparam \mem~67 .shared_arith = "off";

dffeas \mem[6][47] (
	.clk(clk),
	.d(\mem~67_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][47]~q ),
	.prn(vcc));
defparam \mem[6][47] .is_wysiwyg = "true";
defparam \mem[6][47] .power_up = "low";

dffeas \mem[5][47] (
	.clk(clk),
	.d(ShiftLeft147),
	.asdata(\mem[6][47]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][47]~q ),
	.prn(vcc));
defparam \mem[5][47] .is_wysiwyg = "true";
defparam \mem[5][47] .power_up = "low";

dffeas \mem[4][47] (
	.clk(clk),
	.d(ShiftLeft147),
	.asdata(\mem[5][47]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][47]~q ),
	.prn(vcc));
defparam \mem[4][47] .is_wysiwyg = "true";
defparam \mem[4][47] .power_up = "low";

dffeas \mem[3][47] (
	.clk(clk),
	.d(ShiftLeft147),
	.asdata(\mem[4][47]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][47]~q ),
	.prn(vcc));
defparam \mem[3][47] .is_wysiwyg = "true";
defparam \mem[3][47] .power_up = "low";

dffeas \mem[2][47] (
	.clk(clk),
	.d(ShiftLeft147),
	.asdata(\mem[3][47]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][47]~q ),
	.prn(vcc));
defparam \mem[2][47] .is_wysiwyg = "true";
defparam \mem[2][47] .power_up = "low";

dffeas \mem[1][47] (
	.clk(clk),
	.d(ShiftLeft147),
	.asdata(\mem[2][47]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][47]~q ),
	.prn(vcc));
defparam \mem[1][47] .is_wysiwyg = "true";
defparam \mem[1][47] .power_up = "low";

dffeas \mem[7][23] (
	.clk(clk),
	.d(\mem~68_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][23]~q ),
	.prn(vcc));
defparam \mem[7][23] .is_wysiwyg = "true";
defparam \mem[7][23] .power_up = "low";

cyclonev_lcell_comb \mem~68 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft123),
	.datac(!\mem[7][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~68 .extended_lut = "off";
defparam \mem~68 .lut_mask = 64'h2727272727272727;
defparam \mem~68 .shared_arith = "off";

dffeas \mem[6][23] (
	.clk(clk),
	.d(\mem~68_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][23]~q ),
	.prn(vcc));
defparam \mem[6][23] .is_wysiwyg = "true";
defparam \mem[6][23] .power_up = "low";

dffeas \mem[5][23] (
	.clk(clk),
	.d(ShiftLeft123),
	.asdata(\mem[6][23]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][23]~q ),
	.prn(vcc));
defparam \mem[5][23] .is_wysiwyg = "true";
defparam \mem[5][23] .power_up = "low";

dffeas \mem[4][23] (
	.clk(clk),
	.d(ShiftLeft123),
	.asdata(\mem[5][23]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][23]~q ),
	.prn(vcc));
defparam \mem[4][23] .is_wysiwyg = "true";
defparam \mem[4][23] .power_up = "low";

dffeas \mem[3][23] (
	.clk(clk),
	.d(ShiftLeft123),
	.asdata(\mem[4][23]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][23]~q ),
	.prn(vcc));
defparam \mem[3][23] .is_wysiwyg = "true";
defparam \mem[3][23] .power_up = "low";

dffeas \mem[2][23] (
	.clk(clk),
	.d(ShiftLeft123),
	.asdata(\mem[3][23]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][23]~q ),
	.prn(vcc));
defparam \mem[2][23] .is_wysiwyg = "true";
defparam \mem[2][23] .power_up = "low";

dffeas \mem[1][23] (
	.clk(clk),
	.d(ShiftLeft123),
	.asdata(\mem[2][23]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

dffeas \mem[7][55] (
	.clk(clk),
	.d(\mem~69_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][55]~q ),
	.prn(vcc));
defparam \mem[7][55] .is_wysiwyg = "true";
defparam \mem[7][55] .power_up = "low";

cyclonev_lcell_comb \mem~69 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft155),
	.datac(!\mem[7][55]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~69 .extended_lut = "off";
defparam \mem~69 .lut_mask = 64'h2727272727272727;
defparam \mem~69 .shared_arith = "off";

dffeas \mem[6][55] (
	.clk(clk),
	.d(\mem~69_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][55]~q ),
	.prn(vcc));
defparam \mem[6][55] .is_wysiwyg = "true";
defparam \mem[6][55] .power_up = "low";

dffeas \mem[5][55] (
	.clk(clk),
	.d(ShiftLeft155),
	.asdata(\mem[6][55]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][55]~q ),
	.prn(vcc));
defparam \mem[5][55] .is_wysiwyg = "true";
defparam \mem[5][55] .power_up = "low";

dffeas \mem[4][55] (
	.clk(clk),
	.d(ShiftLeft155),
	.asdata(\mem[5][55]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][55]~q ),
	.prn(vcc));
defparam \mem[4][55] .is_wysiwyg = "true";
defparam \mem[4][55] .power_up = "low";

dffeas \mem[3][55] (
	.clk(clk),
	.d(ShiftLeft155),
	.asdata(\mem[4][55]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][55]~q ),
	.prn(vcc));
defparam \mem[3][55] .is_wysiwyg = "true";
defparam \mem[3][55] .power_up = "low";

dffeas \mem[2][55] (
	.clk(clk),
	.d(ShiftLeft155),
	.asdata(\mem[3][55]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][55]~q ),
	.prn(vcc));
defparam \mem[2][55] .is_wysiwyg = "true";
defparam \mem[2][55] .power_up = "low";

dffeas \mem[1][55] (
	.clk(clk),
	.d(ShiftLeft155),
	.asdata(\mem[2][55]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][55]~q ),
	.prn(vcc));
defparam \mem[1][55] .is_wysiwyg = "true";
defparam \mem[1][55] .power_up = "low";

dffeas \mem[7][31] (
	.clk(clk),
	.d(\mem~70_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][31]~q ),
	.prn(vcc));
defparam \mem[7][31] .is_wysiwyg = "true";
defparam \mem[7][31] .power_up = "low";

cyclonev_lcell_comb \mem~70 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft131),
	.datac(!\mem[7][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~70 .extended_lut = "off";
defparam \mem~70 .lut_mask = 64'h2727272727272727;
defparam \mem~70 .shared_arith = "off";

dffeas \mem[6][31] (
	.clk(clk),
	.d(\mem~70_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][31]~q ),
	.prn(vcc));
defparam \mem[6][31] .is_wysiwyg = "true";
defparam \mem[6][31] .power_up = "low";

dffeas \mem[5][31] (
	.clk(clk),
	.d(ShiftLeft131),
	.asdata(\mem[6][31]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][31]~q ),
	.prn(vcc));
defparam \mem[5][31] .is_wysiwyg = "true";
defparam \mem[5][31] .power_up = "low";

dffeas \mem[4][31] (
	.clk(clk),
	.d(ShiftLeft131),
	.asdata(\mem[5][31]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][31]~q ),
	.prn(vcc));
defparam \mem[4][31] .is_wysiwyg = "true";
defparam \mem[4][31] .power_up = "low";

dffeas \mem[3][31] (
	.clk(clk),
	.d(ShiftLeft131),
	.asdata(\mem[4][31]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][31]~q ),
	.prn(vcc));
defparam \mem[3][31] .is_wysiwyg = "true";
defparam \mem[3][31] .power_up = "low";

dffeas \mem[2][31] (
	.clk(clk),
	.d(ShiftLeft131),
	.asdata(\mem[3][31]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][31]~q ),
	.prn(vcc));
defparam \mem[2][31] .is_wysiwyg = "true";
defparam \mem[2][31] .power_up = "low";

dffeas \mem[1][31] (
	.clk(clk),
	.d(ShiftLeft131),
	.asdata(\mem[2][31]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

dffeas \mem[7][63] (
	.clk(clk),
	.d(\mem~71_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][63]~q ),
	.prn(vcc));
defparam \mem[7][63] .is_wysiwyg = "true";
defparam \mem[7][63] .power_up = "low";

cyclonev_lcell_comb \mem~71 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft163),
	.datac(!\mem[7][63]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~71 .extended_lut = "off";
defparam \mem~71 .lut_mask = 64'h2727272727272727;
defparam \mem~71 .shared_arith = "off";

dffeas \mem[6][63] (
	.clk(clk),
	.d(\mem~71_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][63]~q ),
	.prn(vcc));
defparam \mem[6][63] .is_wysiwyg = "true";
defparam \mem[6][63] .power_up = "low";

dffeas \mem[5][63] (
	.clk(clk),
	.d(ShiftLeft163),
	.asdata(\mem[6][63]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][63]~q ),
	.prn(vcc));
defparam \mem[5][63] .is_wysiwyg = "true";
defparam \mem[5][63] .power_up = "low";

dffeas \mem[4][63] (
	.clk(clk),
	.d(ShiftLeft163),
	.asdata(\mem[5][63]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][63]~q ),
	.prn(vcc));
defparam \mem[4][63] .is_wysiwyg = "true";
defparam \mem[4][63] .power_up = "low";

dffeas \mem[3][63] (
	.clk(clk),
	.d(ShiftLeft163),
	.asdata(\mem[4][63]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][63]~q ),
	.prn(vcc));
defparam \mem[3][63] .is_wysiwyg = "true";
defparam \mem[3][63] .power_up = "low";

dffeas \mem[2][63] (
	.clk(clk),
	.d(ShiftLeft163),
	.asdata(\mem[3][63]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][63]~q ),
	.prn(vcc));
defparam \mem[2][63] .is_wysiwyg = "true";
defparam \mem[2][63] .power_up = "low";

dffeas \mem[1][63] (
	.clk(clk),
	.d(ShiftLeft163),
	.asdata(\mem[2][63]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][63]~q ),
	.prn(vcc));
defparam \mem[1][63] .is_wysiwyg = "true";
defparam \mem[1][63] .power_up = "low";

dffeas \mem[7][7] (
	.clk(clk),
	.d(\mem~72_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][7]~q ),
	.prn(vcc));
defparam \mem[7][7] .is_wysiwyg = "true";
defparam \mem[7][7] .power_up = "low";

cyclonev_lcell_comb \mem~72 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft17),
	.datac(!\mem[7][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~72 .extended_lut = "off";
defparam \mem~72 .lut_mask = 64'h2727272727272727;
defparam \mem~72 .shared_arith = "off";

dffeas \mem[6][7] (
	.clk(clk),
	.d(\mem~72_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][7]~q ),
	.prn(vcc));
defparam \mem[6][7] .is_wysiwyg = "true";
defparam \mem[6][7] .power_up = "low";

dffeas \mem[5][7] (
	.clk(clk),
	.d(ShiftLeft17),
	.asdata(\mem[6][7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][7]~q ),
	.prn(vcc));
defparam \mem[5][7] .is_wysiwyg = "true";
defparam \mem[5][7] .power_up = "low";

dffeas \mem[4][7] (
	.clk(clk),
	.d(ShiftLeft17),
	.asdata(\mem[5][7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][7]~q ),
	.prn(vcc));
defparam \mem[4][7] .is_wysiwyg = "true";
defparam \mem[4][7] .power_up = "low";

dffeas \mem[3][7] (
	.clk(clk),
	.d(ShiftLeft17),
	.asdata(\mem[4][7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][7]~q ),
	.prn(vcc));
defparam \mem[3][7] .is_wysiwyg = "true";
defparam \mem[3][7] .power_up = "low";

dffeas \mem[2][7] (
	.clk(clk),
	.d(ShiftLeft17),
	.asdata(\mem[3][7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][7]~q ),
	.prn(vcc));
defparam \mem[2][7] .is_wysiwyg = "true";
defparam \mem[2][7] .power_up = "low";

dffeas \mem[1][7] (
	.clk(clk),
	.d(ShiftLeft17),
	.asdata(\mem[2][7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

dffeas \mem[7][39] (
	.clk(clk),
	.d(\mem~73_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[7][39]~q ),
	.prn(vcc));
defparam \mem[7][39] .is_wysiwyg = "true";
defparam \mem[7][39] .power_up = "low";

cyclonev_lcell_comb \mem~73 (
	.dataa(!mem_used_7),
	.datab(!ShiftLeft139),
	.datac(!\mem[7][39]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~73 .extended_lut = "off";
defparam \mem~73 .lut_mask = 64'h2727272727272727;
defparam \mem~73 .shared_arith = "off";

dffeas \mem[6][39] (
	.clk(clk),
	.d(\mem~73_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][39]~q ),
	.prn(vcc));
defparam \mem[6][39] .is_wysiwyg = "true";
defparam \mem[6][39] .power_up = "low";

dffeas \mem[5][39] (
	.clk(clk),
	.d(ShiftLeft139),
	.asdata(\mem[6][39]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[6]~q ),
	.ena(\always5~0_combout ),
	.q(\mem[5][39]~q ),
	.prn(vcc));
defparam \mem[5][39] .is_wysiwyg = "true";
defparam \mem[5][39] .power_up = "low";

dffeas \mem[4][39] (
	.clk(clk),
	.d(ShiftLeft139),
	.asdata(\mem[5][39]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[5]~q ),
	.ena(\always4~0_combout ),
	.q(\mem[4][39]~q ),
	.prn(vcc));
defparam \mem[4][39] .is_wysiwyg = "true";
defparam \mem[4][39] .power_up = "low";

dffeas \mem[3][39] (
	.clk(clk),
	.d(ShiftLeft139),
	.asdata(\mem[4][39]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[4]~q ),
	.ena(\always3~0_combout ),
	.q(\mem[3][39]~q ),
	.prn(vcc));
defparam \mem[3][39] .is_wysiwyg = "true";
defparam \mem[3][39] .power_up = "low";

dffeas \mem[2][39] (
	.clk(clk),
	.d(ShiftLeft139),
	.asdata(\mem[3][39]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[3]~q ),
	.ena(\always2~0_combout ),
	.q(\mem[2][39]~q ),
	.prn(vcc));
defparam \mem[2][39] .is_wysiwyg = "true";
defparam \mem[2][39] .power_up = "low";

dffeas \mem[1][39] (
	.clk(clk),
	.d(ShiftLeft139),
	.asdata(\mem[2][39]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\mem_used[2]~q ),
	.ena(\always1~0_combout ),
	.q(\mem[1][39]~q ),
	.prn(vcc));
defparam \mem[1][39] .is_wysiwyg = "true";
defparam \mem[1][39] .power_up = "low";

cyclonev_lcell_comb \mem_used[7]~0 (
	.dataa(!mem_used_7),
	.datab(!bready),
	.datac(!\write~0_combout ),
	.datad(!\mem_used[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[7]~0 .extended_lut = "off";
defparam \mem_used[7]~0 .lut_mask = 64'h414D414D414D414D;
defparam \mem_used[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!\write~0_combout ),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h2F3F2F3F2F3F2F3F;
defparam \mem_used[0]~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_master_agent (
	f2h_BVALID_0,
	f2h_RVALID_0,
	mem_68_0,
	mem_64_0,
	mem_69_0,
	mem_65_0,
	mem_70_0,
	mem_66_0,
	mem_71_0,
	mem_67_0,
	mem_68_01,
	mem_64_01,
	mem_used_0,
	src0_valid,
	av_readdatavalid,
	av_readdatavalid1,
	av_readdatavalid2,
	av_readdatavalid3,
	av_readdatavalid4)/* synthesis synthesis_greybox=0 */;
input 	f2h_BVALID_0;
input 	f2h_RVALID_0;
input 	mem_68_0;
input 	mem_64_0;
input 	mem_69_0;
input 	mem_65_0;
input 	mem_70_0;
input 	mem_66_0;
input 	mem_71_0;
input 	mem_67_0;
input 	mem_68_01;
input 	mem_64_01;
input 	mem_used_0;
input 	src0_valid;
output 	av_readdatavalid;
output 	av_readdatavalid1;
output 	av_readdatavalid2;
output 	av_readdatavalid3;
output 	av_readdatavalid4;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \av_readdatavalid~0 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_69_0),
	.datad(!mem_65_0),
	.datae(!mem_70_0),
	.dataf(!mem_66_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdatavalid),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdatavalid~0 .extended_lut = "off";
defparam \av_readdatavalid~0 .lut_mask = 64'h8000000000000000;
defparam \av_readdatavalid~0 .shared_arith = "off";

cyclonev_lcell_comb \av_readdatavalid~1 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdatavalid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdatavalid~1 .extended_lut = "off";
defparam \av_readdatavalid~1 .lut_mask = 64'h8888888888888888;
defparam \av_readdatavalid~1 .shared_arith = "off";

cyclonev_lcell_comb \av_readdatavalid~2 (
	.dataa(!f2h_RVALID_0),
	.datab(!mem_68_01),
	.datac(!mem_64_01),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdatavalid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdatavalid~2 .extended_lut = "off";
defparam \av_readdatavalid~2 .lut_mask = 64'h1515151515151515;
defparam \av_readdatavalid~2 .shared_arith = "off";

cyclonev_lcell_comb \av_readdatavalid~3 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!av_readdatavalid),
	.datae(!av_readdatavalid1),
	.dataf(!av_readdatavalid2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdatavalid3),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdatavalid~3 .extended_lut = "off";
defparam \av_readdatavalid~3 .lut_mask = 64'h01010100FFFFFFFF;
defparam \av_readdatavalid~3 .shared_arith = "off";

cyclonev_lcell_comb \av_readdatavalid~4 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!av_readdatavalid),
	.datae(!av_readdatavalid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdatavalid4),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdatavalid~4 .extended_lut = "off";
defparam \av_readdatavalid~4 .lut_mask = 64'h0101010001010100;
defparam \av_readdatavalid~4 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_traffic_limiter_2 (
	f2h_BVALID_0,
	f2h_RVALID_0,
	clk,
	mem_105_0,
	mem_113_0,
	mem_139_0,
	last_channel_1,
	has_pending_responses1,
	mem_used_0,
	WideOr1,
	reset,
	inc_read,
	bready)/* synthesis synthesis_greybox=0 */;
input 	f2h_BVALID_0;
input 	f2h_RVALID_0;
input 	clk;
input 	mem_105_0;
input 	mem_113_0;
input 	mem_139_0;
output 	last_channel_1;
output 	has_pending_responses1;
input 	mem_used_0;
input 	WideOr1;
input 	reset;
input 	inc_read;
input 	bready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \last_channel[1]~0_combout ;
wire \pending_response_count[0]~1_combout ;
wire \pending_response_count[4]~0_combout ;
wire \pending_response_count[0]~q ;
wire \response_sink_accepted~0_combout ;
wire \Add0~3_combout ;
wire \pending_response_count[1]~q ;
wire \Add0~2_combout ;
wire \pending_response_count[2]~q ;
wire \Add0~1_combout ;
wire \pending_response_count[3]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[4]~q ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~1_combout ;


dffeas \last_channel[1] (
	.clk(clk),
	.d(\last_channel[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

cyclonev_lcell_comb \last_channel[1]~0 (
	.dataa(!last_channel_1),
	.datab(!WideOr1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_channel[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_channel[1]~0 .extended_lut = "off";
defparam \last_channel[1]~0 .lut_mask = 64'h7777777777777777;
defparam \last_channel[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[4]~0 (
	.dataa(!f2h_RVALID_0),
	.datab(!mem_105_0),
	.datac(!inc_read),
	.datad(!mem_113_0),
	.datae(!mem_139_0),
	.dataf(!bready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[4]~0 .extended_lut = "off";
defparam \pending_response_count[4]~0 .lut_mask = 64'hF0A5F0A5F0A53C2D;
defparam \pending_response_count[4]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[4]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!mem_105_0),
	.datae(!mem_113_0),
	.dataf(!mem_139_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h0000333305003733;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~3 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(!\response_sink_accepted~0_combout ),
	.datac(!\pending_response_count[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~3 .extended_lut = "off";
defparam \Add0~3 .lut_mask = 64'h6969696969696969;
defparam \Add0~3 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[4]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(!\response_sink_accepted~0_combout ),
	.datac(!\pending_response_count[2]~q ),
	.datad(!\pending_response_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h2D4B2D4B2D4B2D4B;
defparam \Add0~2 .shared_arith = "off";

dffeas \pending_response_count[2] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[4]~0_combout ),
	.q(\pending_response_count[2]~q ),
	.prn(vcc));
defparam \pending_response_count[2] .is_wysiwyg = "true";
defparam \pending_response_count[2] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(!\response_sink_accepted~0_combout ),
	.datac(!\pending_response_count[3]~q ),
	.datad(!\pending_response_count[2]~q ),
	.datae(!\pending_response_count[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h2D0F0F4B2D0F0F4B;
defparam \Add0~1 .shared_arith = "off";

dffeas \pending_response_count[3] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[4]~0_combout ),
	.q(\pending_response_count[3]~q ),
	.prn(vcc));
defparam \pending_response_count[3] .is_wysiwyg = "true";
defparam \pending_response_count[3] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(!\response_sink_accepted~0_combout ),
	.datac(!\pending_response_count[4]~q ),
	.datad(!\pending_response_count[3]~q ),
	.datae(!\pending_response_count[2]~q ),
	.dataf(!\pending_response_count[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h2D0F0F0F0F0F0F4B;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[4] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[4]~0_combout ),
	.q(\pending_response_count[4]~q ),
	.prn(vcc));
defparam \pending_response_count[4] .is_wysiwyg = "true";
defparam \pending_response_count[4] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!\pending_response_count[4]~q ),
	.datab(!\pending_response_count[3]~q ),
	.datac(!\pending_response_count[2]~q ),
	.datad(!\pending_response_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h8000800080008000;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~1 (
	.dataa(!has_pending_responses1),
	.datab(!inc_read),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(!\has_pending_responses~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~1 .extended_lut = "off";
defparam \has_pending_responses~1 .lut_mask = 64'h5555D5545555D554;
defparam \has_pending_responses~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_width_adapter (
	readaddress_2,
	saved_grant_0,
	ShiftLeft0)/* synthesis synthesis_greybox=0 */;
input 	readaddress_2;
input 	saved_grant_0;
output 	ShiftLeft0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h4444444444444444;
defparam \ShiftLeft0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_width_adapter_2 (
	writeaddress_2,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	writeaddress_1,
	writeaddress_0,
	saved_grant_1,
	last_write_collision,
	last_write_data_0,
	control_2,
	control_0,
	src_payload,
	ShiftLeft1,
	last_write_data_1,
	ShiftLeft11,
	last_write_data_2,
	ShiftLeft12,
	last_write_data_3,
	ShiftLeft13,
	last_write_data_4,
	ShiftLeft14,
	last_write_data_5,
	ShiftLeft15,
	last_write_data_6,
	ShiftLeft16,
	last_write_data_7,
	ShiftLeft17,
	write_writedata,
	last_write_data_8,
	ShiftLeft18,
	write_writedata1,
	last_write_data_9,
	ShiftLeft19,
	write_writedata2,
	last_write_data_10,
	ShiftLeft110,
	write_writedata3,
	last_write_data_11,
	ShiftLeft111,
	write_writedata4,
	last_write_data_12,
	ShiftLeft112,
	write_writedata5,
	last_write_data_13,
	ShiftLeft113,
	write_writedata6,
	last_write_data_14,
	ShiftLeft114,
	write_writedata7,
	last_write_data_15,
	ShiftLeft115,
	last_write_data_16,
	ShiftLeft116,
	last_write_data_17,
	ShiftLeft117,
	last_write_data_18,
	ShiftLeft118,
	last_write_data_19,
	ShiftLeft119,
	last_write_data_20,
	ShiftLeft120,
	last_write_data_21,
	ShiftLeft121,
	last_write_data_22,
	ShiftLeft122,
	last_write_data_23,
	ShiftLeft123,
	last_write_data_24,
	ShiftLeft124,
	last_write_data_25,
	ShiftLeft125,
	last_write_data_26,
	ShiftLeft126,
	last_write_data_27,
	ShiftLeft127,
	last_write_data_28,
	ShiftLeft128,
	last_write_data_29,
	ShiftLeft129,
	last_write_data_30,
	ShiftLeft130,
	last_write_data_31,
	ShiftLeft131,
	ShiftLeft132,
	ShiftLeft133,
	ShiftLeft134,
	ShiftLeft135,
	ShiftLeft136,
	ShiftLeft137,
	ShiftLeft138,
	ShiftLeft139,
	ShiftLeft140,
	ShiftLeft141,
	ShiftLeft142,
	ShiftLeft143,
	ShiftLeft144,
	ShiftLeft145,
	ShiftLeft146,
	ShiftLeft147,
	ShiftLeft148,
	ShiftLeft149,
	ShiftLeft150,
	ShiftLeft151,
	ShiftLeft152,
	ShiftLeft153,
	ShiftLeft154,
	ShiftLeft155,
	ShiftLeft156,
	ShiftLeft157,
	ShiftLeft158,
	ShiftLeft159,
	ShiftLeft160,
	ShiftLeft161,
	ShiftLeft162,
	ShiftLeft163,
	ShiftLeft0,
	ShiftLeft01,
	ShiftLeft02,
	ShiftLeft03,
	ShiftLeft04,
	ShiftLeft05,
	ShiftLeft06,
	ShiftLeft07)/* synthesis synthesis_greybox=0 */;
input 	writeaddress_2;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	writeaddress_1;
input 	writeaddress_0;
input 	saved_grant_1;
input 	last_write_collision;
input 	last_write_data_0;
input 	control_2;
input 	control_0;
input 	src_payload;
output 	ShiftLeft1;
input 	last_write_data_1;
output 	ShiftLeft11;
input 	last_write_data_2;
output 	ShiftLeft12;
input 	last_write_data_3;
output 	ShiftLeft13;
input 	last_write_data_4;
output 	ShiftLeft14;
input 	last_write_data_5;
output 	ShiftLeft15;
input 	last_write_data_6;
output 	ShiftLeft16;
input 	last_write_data_7;
output 	ShiftLeft17;
input 	write_writedata;
input 	last_write_data_8;
output 	ShiftLeft18;
input 	write_writedata1;
input 	last_write_data_9;
output 	ShiftLeft19;
input 	write_writedata2;
input 	last_write_data_10;
output 	ShiftLeft110;
input 	write_writedata3;
input 	last_write_data_11;
output 	ShiftLeft111;
input 	write_writedata4;
input 	last_write_data_12;
output 	ShiftLeft112;
input 	write_writedata5;
input 	last_write_data_13;
output 	ShiftLeft113;
input 	write_writedata6;
input 	last_write_data_14;
output 	ShiftLeft114;
input 	write_writedata7;
input 	last_write_data_15;
output 	ShiftLeft115;
input 	last_write_data_16;
output 	ShiftLeft116;
input 	last_write_data_17;
output 	ShiftLeft117;
input 	last_write_data_18;
output 	ShiftLeft118;
input 	last_write_data_19;
output 	ShiftLeft119;
input 	last_write_data_20;
output 	ShiftLeft120;
input 	last_write_data_21;
output 	ShiftLeft121;
input 	last_write_data_22;
output 	ShiftLeft122;
input 	last_write_data_23;
output 	ShiftLeft123;
input 	last_write_data_24;
output 	ShiftLeft124;
input 	last_write_data_25;
output 	ShiftLeft125;
input 	last_write_data_26;
output 	ShiftLeft126;
input 	last_write_data_27;
output 	ShiftLeft127;
input 	last_write_data_28;
output 	ShiftLeft128;
input 	last_write_data_29;
output 	ShiftLeft129;
input 	last_write_data_30;
output 	ShiftLeft130;
input 	last_write_data_31;
output 	ShiftLeft131;
output 	ShiftLeft132;
output 	ShiftLeft133;
output 	ShiftLeft134;
output 	ShiftLeft135;
output 	ShiftLeft136;
output 	ShiftLeft137;
output 	ShiftLeft138;
output 	ShiftLeft139;
output 	ShiftLeft140;
output 	ShiftLeft141;
output 	ShiftLeft142;
output 	ShiftLeft143;
output 	ShiftLeft144;
output 	ShiftLeft145;
output 	ShiftLeft146;
output 	ShiftLeft147;
output 	ShiftLeft148;
output 	ShiftLeft149;
output 	ShiftLeft150;
output 	ShiftLeft151;
output 	ShiftLeft152;
output 	ShiftLeft153;
output 	ShiftLeft154;
output 	ShiftLeft155;
output 	ShiftLeft156;
output 	ShiftLeft157;
output 	ShiftLeft158;
output 	ShiftLeft159;
output 	ShiftLeft160;
output 	ShiftLeft161;
output 	ShiftLeft162;
output 	ShiftLeft163;
output 	ShiftLeft0;
output 	ShiftLeft01;
output 	ShiftLeft02;
output 	ShiftLeft03;
output 	ShiftLeft04;
output 	ShiftLeft05;
output 	ShiftLeft06;
output 	ShiftLeft07;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ShiftLeft1~8_combout ;
wire \ShiftLeft1~10_combout ;
wire \ShiftLeft1~12_combout ;
wire \ShiftLeft1~14_combout ;
wire \ShiftLeft1~16_combout ;
wire \ShiftLeft1~18_combout ;
wire \ShiftLeft1~20_combout ;
wire \ShiftLeft1~22_combout ;
wire \ShiftLeft1~24_combout ;
wire \ShiftLeft1~26_combout ;
wire \ShiftLeft1~28_combout ;
wire \ShiftLeft1~30_combout ;
wire \ShiftLeft1~32_combout ;
wire \ShiftLeft1~34_combout ;
wire \ShiftLeft1~36_combout ;
wire \ShiftLeft1~38_combout ;
wire \ShiftLeft1~40_combout ;
wire \ShiftLeft1~42_combout ;
wire \ShiftLeft1~44_combout ;
wire \ShiftLeft1~46_combout ;
wire \ShiftLeft1~48_combout ;
wire \ShiftLeft1~50_combout ;
wire \ShiftLeft1~52_combout ;
wire \ShiftLeft1~54_combout ;


cyclonev_lcell_comb \ShiftLeft1~0 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!last_write_data_0),
	.datae(!q_b_0),
	.dataf(!src_payload),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft1),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~0 .extended_lut = "off";
defparam \ShiftLeft1~0 .lut_mask = 64'h00000000000EE0EE;
defparam \ShiftLeft1~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~1 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_1),
	.dataf(!q_b_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft11),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~1 .extended_lut = "off";
defparam \ShiftLeft1~1 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~2 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_2),
	.dataf(!q_b_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft12),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~2 .extended_lut = "off";
defparam \ShiftLeft1~2 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~2 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~3 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_3),
	.dataf(!q_b_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft13),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~3 .extended_lut = "off";
defparam \ShiftLeft1~3 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~4 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_4),
	.dataf(!q_b_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft14),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~4 .extended_lut = "off";
defparam \ShiftLeft1~4 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~4 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~5 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_5),
	.dataf(!q_b_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft15),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~5 .extended_lut = "off";
defparam \ShiftLeft1~5 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~5 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~6 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_6),
	.dataf(!q_b_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft16),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~6 .extended_lut = "off";
defparam \ShiftLeft1~6 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~6 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~7 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_7),
	.dataf(!q_b_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft17),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~7 .extended_lut = "off";
defparam \ShiftLeft1~7 .lut_mask = 64'h0000000E00E000EE;
defparam \ShiftLeft1~7 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~9 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata),
	.datad(!\ShiftLeft1~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft18),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~9 .extended_lut = "off";
defparam \ShiftLeft1~9 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~9 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~11 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata1),
	.datad(!\ShiftLeft1~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft19),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~11 .extended_lut = "off";
defparam \ShiftLeft1~11 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~11 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~13 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata2),
	.datad(!\ShiftLeft1~12_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft110),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~13 .extended_lut = "off";
defparam \ShiftLeft1~13 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~13 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~15 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata3),
	.datad(!\ShiftLeft1~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft111),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~15 .extended_lut = "off";
defparam \ShiftLeft1~15 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~15 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~17 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata4),
	.datad(!\ShiftLeft1~16_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft112),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~17 .extended_lut = "off";
defparam \ShiftLeft1~17 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~17 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~19 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata5),
	.datad(!\ShiftLeft1~18_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft113),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~19 .extended_lut = "off";
defparam \ShiftLeft1~19 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~19 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~21 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata6),
	.datad(!\ShiftLeft1~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft114),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~21 .extended_lut = "off";
defparam \ShiftLeft1~21 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~21 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~23 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata7),
	.datad(!\ShiftLeft1~22_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft115),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~23 .extended_lut = "off";
defparam \ShiftLeft1~23 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~23 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~25 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata),
	.datad(!\ShiftLeft1~24_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft116),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~25 .extended_lut = "off";
defparam \ShiftLeft1~25 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~25 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~27 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata1),
	.datad(!\ShiftLeft1~26_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft117),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~27 .extended_lut = "off";
defparam \ShiftLeft1~27 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~27 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~29 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata2),
	.datad(!\ShiftLeft1~28_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft118),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~29 .extended_lut = "off";
defparam \ShiftLeft1~29 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~29 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~31 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata3),
	.datad(!\ShiftLeft1~30_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft119),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~31 .extended_lut = "off";
defparam \ShiftLeft1~31 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~31 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~33 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata4),
	.datad(!\ShiftLeft1~32_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft120),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~33 .extended_lut = "off";
defparam \ShiftLeft1~33 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~33 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~35 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata5),
	.datad(!\ShiftLeft1~34_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft121),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~35 .extended_lut = "off";
defparam \ShiftLeft1~35 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~35 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~37 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata6),
	.datad(!\ShiftLeft1~36_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft122),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~37 .extended_lut = "off";
defparam \ShiftLeft1~37 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~37 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~39 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata7),
	.datad(!\ShiftLeft1~38_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft123),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~39 .extended_lut = "off";
defparam \ShiftLeft1~39 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~39 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~41 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata),
	.datad(!\ShiftLeft1~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft124),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~41 .extended_lut = "off";
defparam \ShiftLeft1~41 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~41 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~43 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata1),
	.datad(!\ShiftLeft1~42_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft125),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~43 .extended_lut = "off";
defparam \ShiftLeft1~43 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~43 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~45 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata2),
	.datad(!\ShiftLeft1~44_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft126),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~45 .extended_lut = "off";
defparam \ShiftLeft1~45 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~45 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~47 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata3),
	.datad(!\ShiftLeft1~46_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft127),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~47 .extended_lut = "off";
defparam \ShiftLeft1~47 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~47 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~49 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata4),
	.datad(!\ShiftLeft1~48_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft128),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~49 .extended_lut = "off";
defparam \ShiftLeft1~49 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~49 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~51 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata5),
	.datad(!\ShiftLeft1~50_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft129),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~51 .extended_lut = "off";
defparam \ShiftLeft1~51 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~51 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~53 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata6),
	.datad(!\ShiftLeft1~52_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft130),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~53 .extended_lut = "off";
defparam \ShiftLeft1~53 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~53 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~55 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata7),
	.datad(!\ShiftLeft1~54_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft131),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~55 .extended_lut = "off";
defparam \ShiftLeft1~55 .lut_mask = 64'h0444044404440444;
defparam \ShiftLeft1~55 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~56 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!last_write_data_0),
	.datae(!q_b_0),
	.dataf(!src_payload),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft132),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~56 .extended_lut = "off";
defparam \ShiftLeft1~56 .lut_mask = 64'h0000000000011011;
defparam \ShiftLeft1~56 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~57 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_1),
	.dataf(!q_b_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft133),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~57 .extended_lut = "off";
defparam \ShiftLeft1~57 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~57 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~58 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_2),
	.dataf(!q_b_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft134),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~58 .extended_lut = "off";
defparam \ShiftLeft1~58 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~58 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~59 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_3),
	.dataf(!q_b_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft135),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~59 .extended_lut = "off";
defparam \ShiftLeft1~59 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~59 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~60 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_4),
	.dataf(!q_b_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft136),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~60 .extended_lut = "off";
defparam \ShiftLeft1~60 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~60 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~61 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_5),
	.dataf(!q_b_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft137),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~61 .extended_lut = "off";
defparam \ShiftLeft1~61 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~61 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~62 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_6),
	.dataf(!q_b_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft138),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~62 .extended_lut = "off";
defparam \ShiftLeft1~62 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~62 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~63 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!last_write_collision),
	.datad(!src_payload),
	.datae(!last_write_data_7),
	.dataf(!q_b_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft139),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~63 .extended_lut = "off";
defparam \ShiftLeft1~63 .lut_mask = 64'h0000000100100011;
defparam \ShiftLeft1~63 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~64 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata),
	.datad(!\ShiftLeft1~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft140),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~64 .extended_lut = "off";
defparam \ShiftLeft1~64 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~64 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~65 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata1),
	.datad(!\ShiftLeft1~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft141),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~65 .extended_lut = "off";
defparam \ShiftLeft1~65 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~65 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~66 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata2),
	.datad(!\ShiftLeft1~12_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft142),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~66 .extended_lut = "off";
defparam \ShiftLeft1~66 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~66 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~67 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata3),
	.datad(!\ShiftLeft1~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft143),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~67 .extended_lut = "off";
defparam \ShiftLeft1~67 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~67 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~68 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata4),
	.datad(!\ShiftLeft1~16_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft144),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~68 .extended_lut = "off";
defparam \ShiftLeft1~68 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~68 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~69 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata5),
	.datad(!\ShiftLeft1~18_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft145),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~69 .extended_lut = "off";
defparam \ShiftLeft1~69 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~69 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~70 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata6),
	.datad(!\ShiftLeft1~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft146),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~70 .extended_lut = "off";
defparam \ShiftLeft1~70 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~70 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~71 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata7),
	.datad(!\ShiftLeft1~22_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft147),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~71 .extended_lut = "off";
defparam \ShiftLeft1~71 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~71 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~72 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata),
	.datad(!\ShiftLeft1~24_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft148),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~72 .extended_lut = "off";
defparam \ShiftLeft1~72 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~72 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~73 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata1),
	.datad(!\ShiftLeft1~26_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft149),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~73 .extended_lut = "off";
defparam \ShiftLeft1~73 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~73 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~74 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata2),
	.datad(!\ShiftLeft1~28_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft150),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~74 .extended_lut = "off";
defparam \ShiftLeft1~74 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~74 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~75 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata3),
	.datad(!\ShiftLeft1~30_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft151),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~75 .extended_lut = "off";
defparam \ShiftLeft1~75 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~75 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~76 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata4),
	.datad(!\ShiftLeft1~32_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft152),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~76 .extended_lut = "off";
defparam \ShiftLeft1~76 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~76 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~77 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata5),
	.datad(!\ShiftLeft1~34_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft153),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~77 .extended_lut = "off";
defparam \ShiftLeft1~77 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~77 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~78 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata6),
	.datad(!\ShiftLeft1~36_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft154),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~78 .extended_lut = "off";
defparam \ShiftLeft1~78 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~78 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~79 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata7),
	.datad(!\ShiftLeft1~38_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft155),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~79 .extended_lut = "off";
defparam \ShiftLeft1~79 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~79 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~80 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata),
	.datad(!\ShiftLeft1~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft156),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~80 .extended_lut = "off";
defparam \ShiftLeft1~80 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~80 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~81 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata1),
	.datad(!\ShiftLeft1~42_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft157),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~81 .extended_lut = "off";
defparam \ShiftLeft1~81 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~81 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~82 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata2),
	.datad(!\ShiftLeft1~44_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft158),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~82 .extended_lut = "off";
defparam \ShiftLeft1~82 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~82 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~83 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata3),
	.datad(!\ShiftLeft1~46_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft159),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~83 .extended_lut = "off";
defparam \ShiftLeft1~83 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~83 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~84 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata4),
	.datad(!\ShiftLeft1~48_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft160),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~84 .extended_lut = "off";
defparam \ShiftLeft1~84 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~84 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~85 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata5),
	.datad(!\ShiftLeft1~50_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft161),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~85 .extended_lut = "off";
defparam \ShiftLeft1~85 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~85 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~86 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata6),
	.datad(!\ShiftLeft1~52_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft162),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~86 .extended_lut = "off";
defparam \ShiftLeft1~86 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~86 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~87 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!write_writedata7),
	.datad(!\ShiftLeft1~54_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft163),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~87 .extended_lut = "off";
defparam \ShiftLeft1~87 .lut_mask = 64'h0111011101110111;
defparam \ShiftLeft1~87 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h4044404040404040;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft01),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h4040404040444040;
defparam \ShiftLeft0~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft02),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h4040404440404040;
defparam \ShiftLeft0~2 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft03),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h4040404040404044;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft04),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h1011101010101010;
defparam \ShiftLeft0~4 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft05),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "off";
defparam \ShiftLeft0~5 .lut_mask = 64'h1010101010111010;
defparam \ShiftLeft0~5 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~6 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft06),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~6 .extended_lut = "off";
defparam \ShiftLeft0~6 .lut_mask = 64'h1010101110101010;
defparam \ShiftLeft0~6 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~7 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft07),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~7 .extended_lut = "off";
defparam \ShiftLeft0~7 .lut_mask = 64'h1010101010101011;
defparam \ShiftLeft0~7 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~8 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_8),
	.datad(!q_b_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~8 .extended_lut = "off";
defparam \ShiftLeft1~8 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~8 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~10 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_9),
	.datad(!q_b_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~10 .extended_lut = "off";
defparam \ShiftLeft1~10 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~10 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~12 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_10),
	.datad(!q_b_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~12 .extended_lut = "off";
defparam \ShiftLeft1~12 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~12 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~14 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_11),
	.datad(!q_b_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~14 .extended_lut = "off";
defparam \ShiftLeft1~14 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~14 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~16 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_12),
	.datad(!q_b_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~16 .extended_lut = "off";
defparam \ShiftLeft1~16 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~16 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~18 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_13),
	.datad(!q_b_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~18 .extended_lut = "off";
defparam \ShiftLeft1~18 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~18 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~20 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_14),
	.datad(!q_b_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~20 .extended_lut = "off";
defparam \ShiftLeft1~20 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~20 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~22 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_15),
	.datad(!q_b_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~22 .extended_lut = "off";
defparam \ShiftLeft1~22 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~22 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~24 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_16),
	.datad(!q_b_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~24 .extended_lut = "off";
defparam \ShiftLeft1~24 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~24 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~26 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_17),
	.datad(!q_b_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~26 .extended_lut = "off";
defparam \ShiftLeft1~26 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~26 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~28 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_18),
	.datad(!q_b_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~28 .extended_lut = "off";
defparam \ShiftLeft1~28 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~28 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~30 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_19),
	.datad(!q_b_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~30 .extended_lut = "off";
defparam \ShiftLeft1~30 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~30 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~32 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_20),
	.datad(!q_b_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~32 .extended_lut = "off";
defparam \ShiftLeft1~32 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~32 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~34 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_21),
	.datad(!q_b_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~34 .extended_lut = "off";
defparam \ShiftLeft1~34 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~34 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~36 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_22),
	.datad(!q_b_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~36 .extended_lut = "off";
defparam \ShiftLeft1~36 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~36 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~38 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_23),
	.datad(!q_b_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~38 .extended_lut = "off";
defparam \ShiftLeft1~38 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~38 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~40 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_24),
	.datad(!q_b_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~40 .extended_lut = "off";
defparam \ShiftLeft1~40 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~40 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~42 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_25),
	.datad(!q_b_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~42 .extended_lut = "off";
defparam \ShiftLeft1~42 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~42 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~44 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_26),
	.datad(!q_b_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~44 .extended_lut = "off";
defparam \ShiftLeft1~44 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~44 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~46 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_27),
	.datad(!q_b_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~46 .extended_lut = "off";
defparam \ShiftLeft1~46 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~46 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~48 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_28),
	.datad(!q_b_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~48 .extended_lut = "off";
defparam \ShiftLeft1~48 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~48 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~50 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_29),
	.datad(!q_b_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~50 .extended_lut = "off";
defparam \ShiftLeft1~50 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~50 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~52 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_30),
	.datad(!q_b_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~52 .extended_lut = "off";
defparam \ShiftLeft1~52 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~52 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~54 (
	.dataa(!last_write_collision),
	.datab(!control_2),
	.datac(!last_write_data_31),
	.datad(!q_b_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft1~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~54 .extended_lut = "off";
defparam \ShiftLeft1~54 .lut_mask = 64'h048C048C048C048C;
defparam \ShiftLeft1~54 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_1_cmd_demux_001_1 (
	f2h_BVALID_0,
	mem_105_0,
	mem_139_0,
	mem_used_0,
	src0_valid,
	src0_valid1)/* synthesis synthesis_greybox=0 */;
input 	f2h_BVALID_0;
input 	mem_105_0;
input 	mem_139_0;
input 	mem_used_0;
output 	src0_valid;
output 	src0_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!mem_105_0),
	.datab(!mem_139_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h2222222222222222;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~1 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!mem_105_0),
	.datad(!mem_139_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~1 .extended_lut = "off";
defparam \src0_valid~1 .lut_mask = 64'h0010001000100010;
defparam \src0_valid~1 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_1_cmd_mux (
	outclk_wire_0,
	writeaddress_2,
	writeaddress_3,
	writeaddress_4,
	writeaddress_5,
	writeaddress_6,
	writeaddress_7,
	writeaddress_8,
	writeaddress_9,
	writeaddress_10,
	writeaddress_11,
	writeaddress_12,
	writeaddress_13,
	writeaddress_14,
	writeaddress_15,
	writeaddress_16,
	writeaddress_17,
	writeaddress_18,
	writeaddress_19,
	writeaddress_20,
	writeaddress_21,
	writeaddress_22,
	writeaddress_23,
	writeaddress_24,
	writeaddress_25,
	writeaddress_26,
	writeaddress_27,
	writeaddress_28,
	writeaddress_29,
	writeaddress_30,
	writeaddress_31,
	hold_waitrequest,
	fifo_empty,
	saved_grant_1,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	control_2,
	control_0,
	src_payload30,
	altera_reset_synchronizer_int_chain_out,
	write_cp_ready,
	src_payload31)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	writeaddress_2;
input 	writeaddress_3;
input 	writeaddress_4;
input 	writeaddress_5;
input 	writeaddress_6;
input 	writeaddress_7;
input 	writeaddress_8;
input 	writeaddress_9;
input 	writeaddress_10;
input 	writeaddress_11;
input 	writeaddress_12;
input 	writeaddress_13;
input 	writeaddress_14;
input 	writeaddress_15;
input 	writeaddress_16;
input 	writeaddress_17;
input 	writeaddress_18;
input 	writeaddress_19;
input 	writeaddress_20;
input 	writeaddress_21;
input 	writeaddress_22;
input 	writeaddress_23;
input 	writeaddress_24;
input 	writeaddress_25;
input 	writeaddress_26;
input 	writeaddress_27;
input 	writeaddress_28;
input 	writeaddress_29;
input 	writeaddress_30;
input 	writeaddress_31;
input 	hold_waitrequest;
input 	fifo_empty;
output 	saved_grant_1;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
input 	control_2;
input 	control_0;
output 	src_payload30;
input 	altera_reset_synchronizer_int_chain_out;
input 	write_cp_ready;
output 	src_payload31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;


dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\saved_grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!hold_waitrequest),
	.datab(!fifo_empty),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_1),
	.datab(!writeaddress_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_1),
	.datab(!control_2),
	.datac(!control_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h4545454545454545;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!fifo_empty),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!src_valid),
	.datab(!write_cp_ready),
	.datac(!\packet_in_progress~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h4E4E4E4E4E4E4E4E;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!hold_waitrequest),
	.datab(!fifo_empty),
	.datac(!saved_grant_1),
	.datad(!\packet_in_progress~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h110F110F110F110F;
defparam \saved_grant[1]~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_1_cmd_mux_1 (
	f2h_ARREADY_0,
	outclk_wire_0,
	readaddress_2,
	readaddress_3,
	readaddress_4,
	readaddress_5,
	readaddress_6,
	readaddress_7,
	readaddress_8,
	readaddress_9,
	readaddress_10,
	readaddress_11,
	readaddress_12,
	readaddress_13,
	readaddress_14,
	readaddress_15,
	readaddress_16,
	readaddress_17,
	readaddress_18,
	readaddress_19,
	readaddress_20,
	readaddress_21,
	readaddress_22,
	readaddress_23,
	readaddress_24,
	readaddress_25,
	readaddress_26,
	readaddress_27,
	readaddress_28,
	readaddress_29,
	readaddress_30,
	readaddress_31,
	mem_used_7,
	saved_grant_0,
	last_channel_1,
	has_pending_responses,
	read_select,
	hold_waitrequest,
	write,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	altera_reset_synchronizer_int_chain_out,
	WideOr1)/* synthesis synthesis_greybox=0 */;
input 	f2h_ARREADY_0;
input 	outclk_wire_0;
input 	readaddress_2;
input 	readaddress_3;
input 	readaddress_4;
input 	readaddress_5;
input 	readaddress_6;
input 	readaddress_7;
input 	readaddress_8;
input 	readaddress_9;
input 	readaddress_10;
input 	readaddress_11;
input 	readaddress_12;
input 	readaddress_13;
input 	readaddress_14;
input 	readaddress_15;
input 	readaddress_16;
input 	readaddress_17;
input 	readaddress_18;
input 	readaddress_19;
input 	readaddress_20;
input 	readaddress_21;
input 	readaddress_22;
input 	readaddress_23;
input 	readaddress_24;
input 	readaddress_25;
input 	readaddress_26;
input 	readaddress_27;
input 	readaddress_28;
input 	readaddress_29;
input 	readaddress_30;
input 	readaddress_31;
input 	mem_used_7;
output 	saved_grant_0;
input 	last_channel_1;
input 	has_pending_responses;
input 	read_select;
input 	hold_waitrequest;
input 	write;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
input 	altera_reset_synchronizer_int_chain_out;
output 	WideOr1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \saved_grant[0]~0_combout ;


Computer_System_altera_merlin_arbitrator_4 arb(
	.clk(outclk_wire_0),
	.last_channel_1(last_channel_1),
	.has_pending_responses(has_pending_responses),
	.reset(altera_reset_synchronizer_int_chain_out),
	.update_grant(\update_grant~0_combout ),
	.WideOr1(WideOr1),
	.grant_0(\arb|grant[0]~0_combout ));

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\saved_grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!readaddress_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_select),
	.datab(!hold_waitrequest),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr1),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'h1111111111111111;
defparam \WideOr1~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\update_grant~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!f2h_ARREADY_0),
	.datab(!mem_used_7),
	.datac(!write),
	.datad(!\packet_in_progress~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'h0BFB0BFB0BFB0BFB;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!\update_grant~0_combout ),
	.datac(!\arb|grant[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[0]~0 .extended_lut = "off";
defparam \saved_grant[0]~0 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \saved_grant[0]~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_arbitrator_4 (
	clk,
	last_channel_1,
	has_pending_responses,
	reset,
	update_grant,
	WideOr1,
	grant_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	last_channel_1;
input 	has_pending_responses;
input 	reset;
input 	update_grant;
input 	WideOr1;
output 	grant_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!last_channel_1),
	.datab(!has_pending_responses),
	.datac(!WideOr1),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!\top_priority_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'h0D0D000D0D0D000D;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!last_channel_1),
	.datab(!has_pending_responses),
	.datac(!WideOr1),
	.datad(!update_grant),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h0D000D000D000D00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_1_rsp_mux (
	f2h_BVALID_0,
	f2h_RVALID_0,
	f2h_RDATA_0,
	f2h_RDATA_1,
	f2h_RDATA_2,
	f2h_RDATA_3,
	f2h_RDATA_4,
	f2h_RDATA_5,
	f2h_RDATA_6,
	f2h_RDATA_7,
	f2h_RDATA_8,
	f2h_RDATA_9,
	f2h_RDATA_10,
	f2h_RDATA_11,
	f2h_RDATA_12,
	f2h_RDATA_13,
	f2h_RDATA_14,
	f2h_RDATA_15,
	f2h_RDATA_16,
	f2h_RDATA_17,
	f2h_RDATA_18,
	f2h_RDATA_19,
	f2h_RDATA_20,
	f2h_RDATA_21,
	f2h_RDATA_22,
	f2h_RDATA_23,
	f2h_RDATA_24,
	f2h_RDATA_25,
	f2h_RDATA_26,
	f2h_RDATA_27,
	f2h_RDATA_28,
	f2h_RDATA_29,
	f2h_RDATA_30,
	f2h_RDATA_31,
	f2h_RDATA_32,
	f2h_RDATA_33,
	f2h_RDATA_34,
	f2h_RDATA_35,
	f2h_RDATA_36,
	f2h_RDATA_37,
	f2h_RDATA_38,
	f2h_RDATA_39,
	f2h_RDATA_40,
	f2h_RDATA_41,
	f2h_RDATA_42,
	f2h_RDATA_43,
	f2h_RDATA_44,
	f2h_RDATA_45,
	f2h_RDATA_46,
	f2h_RDATA_47,
	f2h_RDATA_48,
	f2h_RDATA_49,
	f2h_RDATA_50,
	f2h_RDATA_51,
	f2h_RDATA_52,
	f2h_RDATA_53,
	f2h_RDATA_54,
	f2h_RDATA_55,
	f2h_RDATA_56,
	f2h_RDATA_57,
	f2h_RDATA_58,
	f2h_RDATA_59,
	f2h_RDATA_60,
	f2h_RDATA_61,
	f2h_RDATA_62,
	f2h_RDATA_63,
	mem_68_0,
	mem_64_0,
	mem_69_0,
	mem_65_0,
	mem_70_0,
	mem_66_0,
	mem_71_0,
	mem_67_0,
	mem_68_01,
	mem_64_01,
	mem_8_0,
	mem_40_0,
	mem_16_0,
	mem_48_0,
	mem_24_0,
	mem_56_0,
	mem_0_0,
	mem_32_0,
	mem_9_0,
	mem_41_0,
	mem_17_0,
	mem_49_0,
	mem_25_0,
	mem_57_0,
	mem_1_0,
	mem_33_0,
	mem_10_0,
	mem_42_0,
	mem_18_0,
	mem_50_0,
	mem_26_0,
	mem_58_0,
	mem_2_0,
	mem_34_0,
	mem_11_0,
	mem_43_0,
	mem_19_0,
	mem_51_0,
	mem_27_0,
	mem_59_0,
	mem_3_0,
	mem_35_0,
	mem_12_0,
	mem_44_0,
	mem_20_0,
	mem_52_0,
	mem_28_0,
	mem_60_0,
	mem_4_0,
	mem_36_0,
	mem_13_0,
	mem_45_0,
	mem_21_0,
	mem_53_0,
	mem_29_0,
	mem_61_0,
	mem_5_0,
	mem_37_0,
	mem_14_0,
	mem_46_0,
	mem_22_0,
	mem_54_0,
	mem_30_0,
	mem_62_0,
	mem_6_0,
	mem_38_0,
	mem_15_0,
	mem_47_0,
	mem_23_0,
	mem_55_0,
	mem_31_0,
	mem_63_0,
	mem_7_0,
	mem_39_0,
	mem_used_0,
	src0_valid,
	src_data_8,
	src_data_81,
	src_data_16,
	src_data_24,
	src_data_0,
	src_data_01,
	src_data_9,
	src_data_91,
	src_data_17,
	src_data_25,
	src_data_1,
	src_data_11,
	src_data_10,
	src_data_101,
	src_data_18,
	src_data_26,
	src_data_2,
	src_data_21,
	src_data_111,
	src_data_112,
	src_data_19,
	src_data_27,
	src_data_3,
	src_data_31,
	src_data_12,
	src_data_121,
	src_data_20,
	src_data_28,
	src_data_4,
	src_data_41,
	src_data_13,
	src_data_131,
	src_data_211,
	src_data_29,
	src_data_5,
	src_data_51,
	src_data_14,
	src_data_141,
	src_data_22,
	src_data_30,
	src_data_6,
	src_data_61,
	src_data_15,
	src_data_151,
	src_data_23,
	src_data_311,
	src_data_7,
	src_data_71,
	src_data_82,
	src_data_92,
	src_data_102,
	src_data_113,
	src_data_122,
	src_data_132,
	src_data_142,
	src_data_152)/* synthesis synthesis_greybox=0 */;
input 	f2h_BVALID_0;
input 	f2h_RVALID_0;
input 	f2h_RDATA_0;
input 	f2h_RDATA_1;
input 	f2h_RDATA_2;
input 	f2h_RDATA_3;
input 	f2h_RDATA_4;
input 	f2h_RDATA_5;
input 	f2h_RDATA_6;
input 	f2h_RDATA_7;
input 	f2h_RDATA_8;
input 	f2h_RDATA_9;
input 	f2h_RDATA_10;
input 	f2h_RDATA_11;
input 	f2h_RDATA_12;
input 	f2h_RDATA_13;
input 	f2h_RDATA_14;
input 	f2h_RDATA_15;
input 	f2h_RDATA_16;
input 	f2h_RDATA_17;
input 	f2h_RDATA_18;
input 	f2h_RDATA_19;
input 	f2h_RDATA_20;
input 	f2h_RDATA_21;
input 	f2h_RDATA_22;
input 	f2h_RDATA_23;
input 	f2h_RDATA_24;
input 	f2h_RDATA_25;
input 	f2h_RDATA_26;
input 	f2h_RDATA_27;
input 	f2h_RDATA_28;
input 	f2h_RDATA_29;
input 	f2h_RDATA_30;
input 	f2h_RDATA_31;
input 	f2h_RDATA_32;
input 	f2h_RDATA_33;
input 	f2h_RDATA_34;
input 	f2h_RDATA_35;
input 	f2h_RDATA_36;
input 	f2h_RDATA_37;
input 	f2h_RDATA_38;
input 	f2h_RDATA_39;
input 	f2h_RDATA_40;
input 	f2h_RDATA_41;
input 	f2h_RDATA_42;
input 	f2h_RDATA_43;
input 	f2h_RDATA_44;
input 	f2h_RDATA_45;
input 	f2h_RDATA_46;
input 	f2h_RDATA_47;
input 	f2h_RDATA_48;
input 	f2h_RDATA_49;
input 	f2h_RDATA_50;
input 	f2h_RDATA_51;
input 	f2h_RDATA_52;
input 	f2h_RDATA_53;
input 	f2h_RDATA_54;
input 	f2h_RDATA_55;
input 	f2h_RDATA_56;
input 	f2h_RDATA_57;
input 	f2h_RDATA_58;
input 	f2h_RDATA_59;
input 	f2h_RDATA_60;
input 	f2h_RDATA_61;
input 	f2h_RDATA_62;
input 	f2h_RDATA_63;
input 	mem_68_0;
input 	mem_64_0;
input 	mem_69_0;
input 	mem_65_0;
input 	mem_70_0;
input 	mem_66_0;
input 	mem_71_0;
input 	mem_67_0;
input 	mem_68_01;
input 	mem_64_01;
input 	mem_8_0;
input 	mem_40_0;
input 	mem_16_0;
input 	mem_48_0;
input 	mem_24_0;
input 	mem_56_0;
input 	mem_0_0;
input 	mem_32_0;
input 	mem_9_0;
input 	mem_41_0;
input 	mem_17_0;
input 	mem_49_0;
input 	mem_25_0;
input 	mem_57_0;
input 	mem_1_0;
input 	mem_33_0;
input 	mem_10_0;
input 	mem_42_0;
input 	mem_18_0;
input 	mem_50_0;
input 	mem_26_0;
input 	mem_58_0;
input 	mem_2_0;
input 	mem_34_0;
input 	mem_11_0;
input 	mem_43_0;
input 	mem_19_0;
input 	mem_51_0;
input 	mem_27_0;
input 	mem_59_0;
input 	mem_3_0;
input 	mem_35_0;
input 	mem_12_0;
input 	mem_44_0;
input 	mem_20_0;
input 	mem_52_0;
input 	mem_28_0;
input 	mem_60_0;
input 	mem_4_0;
input 	mem_36_0;
input 	mem_13_0;
input 	mem_45_0;
input 	mem_21_0;
input 	mem_53_0;
input 	mem_29_0;
input 	mem_61_0;
input 	mem_5_0;
input 	mem_37_0;
input 	mem_14_0;
input 	mem_46_0;
input 	mem_22_0;
input 	mem_54_0;
input 	mem_30_0;
input 	mem_62_0;
input 	mem_6_0;
input 	mem_38_0;
input 	mem_15_0;
input 	mem_47_0;
input 	mem_23_0;
input 	mem_55_0;
input 	mem_31_0;
input 	mem_63_0;
input 	mem_7_0;
input 	mem_39_0;
input 	mem_used_0;
input 	src0_valid;
output 	src_data_8;
output 	src_data_81;
output 	src_data_16;
output 	src_data_24;
output 	src_data_0;
output 	src_data_01;
output 	src_data_9;
output 	src_data_91;
output 	src_data_17;
output 	src_data_25;
output 	src_data_1;
output 	src_data_11;
output 	src_data_10;
output 	src_data_101;
output 	src_data_18;
output 	src_data_26;
output 	src_data_2;
output 	src_data_21;
output 	src_data_111;
output 	src_data_112;
output 	src_data_19;
output 	src_data_27;
output 	src_data_3;
output 	src_data_31;
output 	src_data_12;
output 	src_data_121;
output 	src_data_20;
output 	src_data_28;
output 	src_data_4;
output 	src_data_41;
output 	src_data_13;
output 	src_data_131;
output 	src_data_211;
output 	src_data_29;
output 	src_data_5;
output 	src_data_51;
output 	src_data_14;
output 	src_data_141;
output 	src_data_22;
output 	src_data_30;
output 	src_data_6;
output 	src_data_61;
output 	src_data_15;
output 	src_data_151;
output 	src_data_23;
output 	src_data_311;
output 	src_data_7;
output 	src_data_71;
output 	src_data_82;
output 	src_data_92;
output 	src_data_102;
output 	src_data_113;
output 	src_data_122;
output 	src_data_132;
output 	src_data_142;
output 	src_data_152;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_data[16]~2_combout ;
wire \src_data[16]~3_combout ;
wire \src_data[24]~5_combout ;
wire \src_data[24]~6_combout ;
wire \src_data[17]~12_combout ;
wire \src_data[17]~13_combout ;
wire \src_data[25]~15_combout ;
wire \src_data[25]~16_combout ;
wire \src_data[18]~22_combout ;
wire \src_data[18]~23_combout ;
wire \src_data[26]~25_combout ;
wire \src_data[26]~26_combout ;
wire \src_data[19]~32_combout ;
wire \src_data[19]~33_combout ;
wire \src_data[27]~35_combout ;
wire \src_data[27]~36_combout ;
wire \src_data[20]~42_combout ;
wire \src_data[20]~43_combout ;
wire \src_data[28]~45_combout ;
wire \src_data[28]~46_combout ;
wire \src_data[21]~52_combout ;
wire \src_data[21]~53_combout ;
wire \src_data[29]~55_combout ;
wire \src_data[29]~56_combout ;
wire \src_data[22]~62_combout ;
wire \src_data[22]~63_combout ;
wire \src_data[30]~65_combout ;
wire \src_data[30]~66_combout ;
wire \src_data[23]~72_combout ;
wire \src_data[23]~73_combout ;
wire \src_data[31]~75_combout ;
wire \src_data[31]~76_combout ;


cyclonev_lcell_comb \src_data[8]~0 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_8_0),
	.datad(!mem_40_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~0 .extended_lut = "off";
defparam \src_data[8]~0 .lut_mask = 64'h0357035703570357;
defparam \src_data[8]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~1 (
	.dataa(!f2h_RDATA_8),
	.datab(!f2h_RDATA_40),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_81),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~1 .extended_lut = "off";
defparam \src_data[8]~1 .lut_mask = 64'h0357035703570357;
defparam \src_data[8]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~4 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[16]~2_combout ),
	.datae(!\src_data[16]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~4 .extended_lut = "off";
defparam \src_data[16]~4 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[16]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~7 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[24]~5_combout ),
	.datae(!\src_data[24]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~7 .extended_lut = "off";
defparam \src_data[24]~7 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[24]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~8 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_0_0),
	.datad(!mem_32_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~8 .extended_lut = "off";
defparam \src_data[0]~8 .lut_mask = 64'h0357035703570357;
defparam \src_data[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~9 (
	.dataa(!f2h_RDATA_0),
	.datab(!f2h_RDATA_32),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~9 .extended_lut = "off";
defparam \src_data[0]~9 .lut_mask = 64'h0357035703570357;
defparam \src_data[0]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~10 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_9_0),
	.datad(!mem_41_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~10 .extended_lut = "off";
defparam \src_data[9]~10 .lut_mask = 64'h0357035703570357;
defparam \src_data[9]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~11 (
	.dataa(!f2h_RDATA_9),
	.datab(!f2h_RDATA_41),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~11 .extended_lut = "off";
defparam \src_data[9]~11 .lut_mask = 64'h0357035703570357;
defparam \src_data[9]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~14 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[17]~12_combout ),
	.datae(!\src_data[17]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~14 .extended_lut = "off";
defparam \src_data[17]~14 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[17]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~17 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[25]~15_combout ),
	.datae(!\src_data[25]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~17 .extended_lut = "off";
defparam \src_data[25]~17 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[25]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~18 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_1_0),
	.datad(!mem_33_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~18 .extended_lut = "off";
defparam \src_data[1]~18 .lut_mask = 64'h0357035703570357;
defparam \src_data[1]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~19 (
	.dataa(!f2h_RDATA_1),
	.datab(!f2h_RDATA_33),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~19 .extended_lut = "off";
defparam \src_data[1]~19 .lut_mask = 64'h0357035703570357;
defparam \src_data[1]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~20 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_10_0),
	.datad(!mem_42_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~20 .extended_lut = "off";
defparam \src_data[10]~20 .lut_mask = 64'h0357035703570357;
defparam \src_data[10]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~21 (
	.dataa(!f2h_RDATA_10),
	.datab(!f2h_RDATA_42),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~21 .extended_lut = "off";
defparam \src_data[10]~21 .lut_mask = 64'h0357035703570357;
defparam \src_data[10]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~24 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[18]~22_combout ),
	.datae(!\src_data[18]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~24 .extended_lut = "off";
defparam \src_data[18]~24 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[18]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~27 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[26]~25_combout ),
	.datae(!\src_data[26]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~27 .extended_lut = "off";
defparam \src_data[26]~27 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[26]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~28 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_2_0),
	.datad(!mem_34_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~28 .extended_lut = "off";
defparam \src_data[2]~28 .lut_mask = 64'h0357035703570357;
defparam \src_data[2]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~29 (
	.dataa(!f2h_RDATA_2),
	.datab(!f2h_RDATA_34),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~29 .extended_lut = "off";
defparam \src_data[2]~29 .lut_mask = 64'h0357035703570357;
defparam \src_data[2]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~30 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_11_0),
	.datad(!mem_43_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~30 .extended_lut = "off";
defparam \src_data[11]~30 .lut_mask = 64'h0357035703570357;
defparam \src_data[11]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~31 (
	.dataa(!f2h_RDATA_11),
	.datab(!f2h_RDATA_43),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~31 .extended_lut = "off";
defparam \src_data[11]~31 .lut_mask = 64'h0357035703570357;
defparam \src_data[11]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~34 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[19]~32_combout ),
	.datae(!\src_data[19]~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~34 .extended_lut = "off";
defparam \src_data[19]~34 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[19]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~37 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[27]~35_combout ),
	.datae(!\src_data[27]~36_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~37 .extended_lut = "off";
defparam \src_data[27]~37 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[27]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~38 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_3_0),
	.datad(!mem_35_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~38 .extended_lut = "off";
defparam \src_data[3]~38 .lut_mask = 64'h0357035703570357;
defparam \src_data[3]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~39 (
	.dataa(!f2h_RDATA_3),
	.datab(!f2h_RDATA_35),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~39 .extended_lut = "off";
defparam \src_data[3]~39 .lut_mask = 64'h0357035703570357;
defparam \src_data[3]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~40 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_12_0),
	.datad(!mem_44_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~40 .extended_lut = "off";
defparam \src_data[12]~40 .lut_mask = 64'h0357035703570357;
defparam \src_data[12]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~41 (
	.dataa(!f2h_RDATA_12),
	.datab(!f2h_RDATA_44),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_121),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~41 .extended_lut = "off";
defparam \src_data[12]~41 .lut_mask = 64'h0357035703570357;
defparam \src_data[12]~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~44 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[20]~42_combout ),
	.datae(!\src_data[20]~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~44 .extended_lut = "off";
defparam \src_data[20]~44 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[20]~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~47 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[28]~45_combout ),
	.datae(!\src_data[28]~46_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~47 .extended_lut = "off";
defparam \src_data[28]~47 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[28]~47 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~48 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_4_0),
	.datad(!mem_36_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~48 .extended_lut = "off";
defparam \src_data[4]~48 .lut_mask = 64'h0357035703570357;
defparam \src_data[4]~48 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~49 (
	.dataa(!f2h_RDATA_4),
	.datab(!f2h_RDATA_36),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~49 .extended_lut = "off";
defparam \src_data[4]~49 .lut_mask = 64'h0357035703570357;
defparam \src_data[4]~49 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~50 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_13_0),
	.datad(!mem_45_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~50 .extended_lut = "off";
defparam \src_data[13]~50 .lut_mask = 64'h0357035703570357;
defparam \src_data[13]~50 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~51 (
	.dataa(!f2h_RDATA_13),
	.datab(!f2h_RDATA_45),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_131),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~51 .extended_lut = "off";
defparam \src_data[13]~51 .lut_mask = 64'h0357035703570357;
defparam \src_data[13]~51 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~54 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[21]~52_combout ),
	.datae(!\src_data[21]~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_211),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~54 .extended_lut = "off";
defparam \src_data[21]~54 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[21]~54 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~57 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[29]~55_combout ),
	.datae(!\src_data[29]~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~57 .extended_lut = "off";
defparam \src_data[29]~57 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[29]~57 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~58 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_5_0),
	.datad(!mem_37_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~58 .extended_lut = "off";
defparam \src_data[5]~58 .lut_mask = 64'h0357035703570357;
defparam \src_data[5]~58 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~59 (
	.dataa(!f2h_RDATA_5),
	.datab(!f2h_RDATA_37),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~59 .extended_lut = "off";
defparam \src_data[5]~59 .lut_mask = 64'h0357035703570357;
defparam \src_data[5]~59 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~60 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_14_0),
	.datad(!mem_46_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~60 .extended_lut = "off";
defparam \src_data[14]~60 .lut_mask = 64'h0357035703570357;
defparam \src_data[14]~60 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~61 (
	.dataa(!f2h_RDATA_14),
	.datab(!f2h_RDATA_46),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_141),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~61 .extended_lut = "off";
defparam \src_data[14]~61 .lut_mask = 64'h0357035703570357;
defparam \src_data[14]~61 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~64 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[22]~62_combout ),
	.datae(!\src_data[22]~63_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~64 .extended_lut = "off";
defparam \src_data[22]~64 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[22]~64 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~67 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[30]~65_combout ),
	.datae(!\src_data[30]~66_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~67 .extended_lut = "off";
defparam \src_data[30]~67 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[30]~67 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~68 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_6_0),
	.datad(!mem_38_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~68 .extended_lut = "off";
defparam \src_data[6]~68 .lut_mask = 64'h0357035703570357;
defparam \src_data[6]~68 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~69 (
	.dataa(!f2h_RDATA_6),
	.datab(!f2h_RDATA_38),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_61),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~69 .extended_lut = "off";
defparam \src_data[6]~69 .lut_mask = 64'h0357035703570357;
defparam \src_data[6]~69 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~70 (
	.dataa(!mem_69_0),
	.datab(!mem_65_0),
	.datac(!mem_15_0),
	.datad(!mem_47_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~70 .extended_lut = "off";
defparam \src_data[15]~70 .lut_mask = 64'h0357035703570357;
defparam \src_data[15]~70 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~71 (
	.dataa(!f2h_RDATA_15),
	.datab(!f2h_RDATA_47),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_151),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~71 .extended_lut = "off";
defparam \src_data[15]~71 .lut_mask = 64'h0357035703570357;
defparam \src_data[15]~71 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~74 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[23]~72_combout ),
	.datae(!\src_data[23]~73_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~74 .extended_lut = "off";
defparam \src_data[23]~74 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[23]~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~77 (
	.dataa(!f2h_BVALID_0),
	.datab(!mem_used_0),
	.datac(!src0_valid),
	.datad(!\src_data[31]~75_combout ),
	.datae(!\src_data[31]~76_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_311),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~77 .extended_lut = "off";
defparam \src_data[31]~77 .lut_mask = 64'h0001FFFF0001FFFF;
defparam \src_data[31]~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~78 (
	.dataa(!mem_68_0),
	.datab(!mem_64_0),
	.datac(!mem_7_0),
	.datad(!mem_39_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~78 .extended_lut = "off";
defparam \src_data[7]~78 .lut_mask = 64'h0357035703570357;
defparam \src_data[7]~78 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~79 (
	.dataa(!f2h_RDATA_7),
	.datab(!f2h_RDATA_39),
	.datac(!mem_68_01),
	.datad(!mem_64_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~79 .extended_lut = "off";
defparam \src_data[7]~79 .lut_mask = 64'h0357035703570357;
defparam \src_data[7]~79 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~80 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_8),
	.dataf(!src_data_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~80 .extended_lut = "off";
defparam \src_data[8]~80 .lut_mask = 64'h0000000533333337;
defparam \src_data[8]~80 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~81 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_9),
	.dataf(!src_data_91),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~81 .extended_lut = "off";
defparam \src_data[9]~81 .lut_mask = 64'h0000000533333337;
defparam \src_data[9]~81 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~82 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_10),
	.dataf(!src_data_101),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~82 .extended_lut = "off";
defparam \src_data[10]~82 .lut_mask = 64'h0000000533333337;
defparam \src_data[10]~82 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~83 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_111),
	.dataf(!src_data_112),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_113),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~83 .extended_lut = "off";
defparam \src_data[11]~83 .lut_mask = 64'h0000000533333337;
defparam \src_data[11]~83 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~84 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_12),
	.dataf(!src_data_121),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_122),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~84 .extended_lut = "off";
defparam \src_data[12]~84 .lut_mask = 64'h0000000533333337;
defparam \src_data[12]~84 .shared_arith = "off";

cyclonev_lcell_comb \src_data[13]~85 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_13),
	.dataf(!src_data_131),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_132),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13]~85 .extended_lut = "off";
defparam \src_data[13]~85 .lut_mask = 64'h0000000533333337;
defparam \src_data[13]~85 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~86 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_14),
	.dataf(!src_data_141),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_142),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~86 .extended_lut = "off";
defparam \src_data[14]~86 .lut_mask = 64'h0000000533333337;
defparam \src_data[14]~86 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~87 (
	.dataa(!f2h_BVALID_0),
	.datab(!f2h_RVALID_0),
	.datac(!mem_used_0),
	.datad(!src0_valid),
	.datae(!src_data_15),
	.dataf(!src_data_151),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_152),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~87 .extended_lut = "off";
defparam \src_data[15]~87 .lut_mask = 64'h0000000533333337;
defparam \src_data[15]~87 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~2 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_16_0),
	.datad(!mem_48_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[16]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~2 .extended_lut = "off";
defparam \src_data[16]~2 .lut_mask = 64'h0357035703570357;
defparam \src_data[16]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~3 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_16),
	.datac(!f2h_RDATA_48),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[16]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~3 .extended_lut = "off";
defparam \src_data[16]~3 .lut_mask = 64'h0005111500051115;
defparam \src_data[16]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~5 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_24_0),
	.datad(!mem_56_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[24]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~5 .extended_lut = "off";
defparam \src_data[24]~5 .lut_mask = 64'h0357035703570357;
defparam \src_data[24]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[24]~6 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_24),
	.datac(!f2h_RDATA_56),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[24]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24]~6 .extended_lut = "off";
defparam \src_data[24]~6 .lut_mask = 64'h0005111500051115;
defparam \src_data[24]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~12 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_17_0),
	.datad(!mem_49_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[17]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~12 .extended_lut = "off";
defparam \src_data[17]~12 .lut_mask = 64'h0357035703570357;
defparam \src_data[17]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[17]~13 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_17),
	.datac(!f2h_RDATA_49),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[17]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17]~13 .extended_lut = "off";
defparam \src_data[17]~13 .lut_mask = 64'h0005111500051115;
defparam \src_data[17]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~15 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_25_0),
	.datad(!mem_57_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[25]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~15 .extended_lut = "off";
defparam \src_data[25]~15 .lut_mask = 64'h0357035703570357;
defparam \src_data[25]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~16 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_25),
	.datac(!f2h_RDATA_57),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[25]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~16 .extended_lut = "off";
defparam \src_data[25]~16 .lut_mask = 64'h0005111500051115;
defparam \src_data[25]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~22 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_18_0),
	.datad(!mem_50_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[18]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~22 .extended_lut = "off";
defparam \src_data[18]~22 .lut_mask = 64'h0357035703570357;
defparam \src_data[18]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~23 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_18),
	.datac(!f2h_RDATA_50),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[18]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~23 .extended_lut = "off";
defparam \src_data[18]~23 .lut_mask = 64'h0005111500051115;
defparam \src_data[18]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~25 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_26_0),
	.datad(!mem_58_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[26]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~25 .extended_lut = "off";
defparam \src_data[26]~25 .lut_mask = 64'h0357035703570357;
defparam \src_data[26]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~26 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_26),
	.datac(!f2h_RDATA_58),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~26 .extended_lut = "off";
defparam \src_data[26]~26 .lut_mask = 64'h0005111500051115;
defparam \src_data[26]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~32 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_19_0),
	.datad(!mem_51_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[19]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~32 .extended_lut = "off";
defparam \src_data[19]~32 .lut_mask = 64'h0357035703570357;
defparam \src_data[19]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~33 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_19),
	.datac(!f2h_RDATA_51),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[19]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~33 .extended_lut = "off";
defparam \src_data[19]~33 .lut_mask = 64'h0005111500051115;
defparam \src_data[19]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~35 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_27_0),
	.datad(!mem_59_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~35 .extended_lut = "off";
defparam \src_data[27]~35 .lut_mask = 64'h0357035703570357;
defparam \src_data[27]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~36 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_27),
	.datac(!f2h_RDATA_59),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~36 .extended_lut = "off";
defparam \src_data[27]~36 .lut_mask = 64'h0005111500051115;
defparam \src_data[27]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~42 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_20_0),
	.datad(!mem_52_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[20]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~42 .extended_lut = "off";
defparam \src_data[20]~42 .lut_mask = 64'h0357035703570357;
defparam \src_data[20]~42 .shared_arith = "off";

cyclonev_lcell_comb \src_data[20]~43 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_20),
	.datac(!f2h_RDATA_52),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[20]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20]~43 .extended_lut = "off";
defparam \src_data[20]~43 .lut_mask = 64'h0005111500051115;
defparam \src_data[20]~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~45 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_28_0),
	.datad(!mem_60_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~45 .extended_lut = "off";
defparam \src_data[28]~45 .lut_mask = 64'h0357035703570357;
defparam \src_data[28]~45 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~46 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_28),
	.datac(!f2h_RDATA_60),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~46 .extended_lut = "off";
defparam \src_data[28]~46 .lut_mask = 64'h0005111500051115;
defparam \src_data[28]~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~52 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_21_0),
	.datad(!mem_53_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[21]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~52 .extended_lut = "off";
defparam \src_data[21]~52 .lut_mask = 64'h0357035703570357;
defparam \src_data[21]~52 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~53 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_21),
	.datac(!f2h_RDATA_53),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[21]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~53 .extended_lut = "off";
defparam \src_data[21]~53 .lut_mask = 64'h0005111500051115;
defparam \src_data[21]~53 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~55 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_29_0),
	.datad(!mem_61_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[29]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~55 .extended_lut = "off";
defparam \src_data[29]~55 .lut_mask = 64'h0357035703570357;
defparam \src_data[29]~55 .shared_arith = "off";

cyclonev_lcell_comb \src_data[29]~56 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_29),
	.datac(!f2h_RDATA_61),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[29]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29]~56 .extended_lut = "off";
defparam \src_data[29]~56 .lut_mask = 64'h0005111500051115;
defparam \src_data[29]~56 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~62 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_22_0),
	.datad(!mem_54_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[22]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~62 .extended_lut = "off";
defparam \src_data[22]~62 .lut_mask = 64'h0357035703570357;
defparam \src_data[22]~62 .shared_arith = "off";

cyclonev_lcell_comb \src_data[22]~63 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_22),
	.datac(!f2h_RDATA_54),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[22]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22]~63 .extended_lut = "off";
defparam \src_data[22]~63 .lut_mask = 64'h0005111500051115;
defparam \src_data[22]~63 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~65 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_30_0),
	.datad(!mem_62_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~65 .extended_lut = "off";
defparam \src_data[30]~65 .lut_mask = 64'h0357035703570357;
defparam \src_data[30]~65 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~66 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_30),
	.datac(!f2h_RDATA_62),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~66 .extended_lut = "off";
defparam \src_data[30]~66 .lut_mask = 64'h0005111500051115;
defparam \src_data[30]~66 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~72 (
	.dataa(!mem_70_0),
	.datab(!mem_66_0),
	.datac(!mem_23_0),
	.datad(!mem_55_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[23]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~72 .extended_lut = "off";
defparam \src_data[23]~72 .lut_mask = 64'h0357035703570357;
defparam \src_data[23]~72 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~73 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_23),
	.datac(!f2h_RDATA_55),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[23]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~73 .extended_lut = "off";
defparam \src_data[23]~73 .lut_mask = 64'h0005111500051115;
defparam \src_data[23]~73 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~75 (
	.dataa(!mem_71_0),
	.datab(!mem_67_0),
	.datac(!mem_31_0),
	.datad(!mem_63_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[31]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~75 .extended_lut = "off";
defparam \src_data[31]~75 .lut_mask = 64'h0357035703570357;
defparam \src_data[31]~75 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~76 (
	.dataa(!f2h_RVALID_0),
	.datab(!f2h_RDATA_31),
	.datac(!f2h_RDATA_63),
	.datad(!mem_68_01),
	.datae(!mem_64_01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[31]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~76 .extended_lut = "off";
defparam \src_data[31]~76 .lut_mask = 64'h0005111500051115;
defparam \src_data[31]~76 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_2 (
	outclk_wire_0,
	readaddress_15,
	writeaddress_15,
	q_b_0,
	readaddress_2,
	writeaddress_2,
	readaddress_3,
	writeaddress_3,
	readaddress_4,
	writeaddress_4,
	readaddress_5,
	writeaddress_5,
	readaddress_6,
	writeaddress_6,
	readaddress_7,
	writeaddress_7,
	readaddress_8,
	writeaddress_8,
	readaddress_9,
	writeaddress_9,
	readaddress_10,
	writeaddress_10,
	readaddress_11,
	writeaddress_11,
	readaddress_12,
	writeaddress_12,
	readaddress_13,
	writeaddress_13,
	readaddress_14,
	writeaddress_14,
	writeaddress_1,
	writeaddress_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	hold_waitrequest,
	saved_grant_0,
	saved_grant_1,
	mem_used_1,
	fifo_empty,
	last_write_collision,
	last_write_data_0,
	control_2,
	control_0,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	last_write_data_1,
	src_payload1,
	last_write_data_2,
	src_payload2,
	last_write_data_3,
	src_payload3,
	last_write_data_4,
	src_payload4,
	last_write_data_5,
	src_payload5,
	last_write_data_6,
	src_payload6,
	last_write_data_7,
	src_payload7,
	write_writedata,
	last_write_data_8,
	src_payload8,
	src_data_33,
	write_writedata1,
	last_write_data_9,
	src_payload9,
	write_writedata2,
	last_write_data_10,
	src_payload10,
	write_writedata3,
	last_write_data_11,
	src_payload11,
	write_writedata4,
	last_write_data_12,
	src_payload12,
	write_writedata5,
	last_write_data_13,
	src_payload13,
	write_writedata6,
	last_write_data_14,
	src_payload14,
	write_writedata7,
	last_write_data_15,
	src_payload15,
	last_write_data_16,
	src_payload16,
	src_data_34,
	last_write_data_17,
	src_payload17,
	last_write_data_18,
	src_payload18,
	last_write_data_19,
	src_payload19,
	last_write_data_20,
	src_payload20,
	last_write_data_21,
	src_payload21,
	last_write_data_22,
	src_payload22,
	last_write_data_23,
	src_payload23,
	last_write_data_24,
	src_payload24,
	src_data_35,
	last_write_data_25,
	src_payload25,
	last_write_data_26,
	src_payload26,
	last_write_data_27,
	src_payload27,
	last_write_data_28,
	src_payload28,
	last_write_data_29,
	src_payload29,
	last_write_data_30,
	src_payload30,
	last_write_data_31,
	src_payload31,
	r_sync_rst,
	src0_valid,
	read_select,
	read_latency_shift_reg,
	src_data_51)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	readaddress_15;
input 	writeaddress_15;
input 	q_b_0;
input 	readaddress_2;
input 	writeaddress_2;
input 	readaddress_3;
input 	writeaddress_3;
input 	readaddress_4;
input 	writeaddress_4;
input 	readaddress_5;
input 	writeaddress_5;
input 	readaddress_6;
input 	writeaddress_6;
input 	readaddress_7;
input 	writeaddress_7;
input 	readaddress_8;
input 	writeaddress_8;
input 	readaddress_9;
input 	writeaddress_9;
input 	readaddress_10;
input 	writeaddress_10;
input 	readaddress_11;
input 	writeaddress_11;
input 	readaddress_12;
input 	writeaddress_12;
input 	readaddress_13;
input 	writeaddress_13;
input 	readaddress_14;
input 	writeaddress_14;
input 	writeaddress_1;
input 	writeaddress_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
output 	hold_waitrequest;
output 	saved_grant_0;
output 	saved_grant_1;
output 	mem_used_1;
input 	fifo_empty;
input 	last_write_collision;
input 	last_write_data_0;
input 	control_2;
input 	control_0;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_32;
input 	last_write_data_1;
output 	src_payload1;
input 	last_write_data_2;
output 	src_payload2;
input 	last_write_data_3;
output 	src_payload3;
input 	last_write_data_4;
output 	src_payload4;
input 	last_write_data_5;
output 	src_payload5;
input 	last_write_data_6;
output 	src_payload6;
input 	last_write_data_7;
output 	src_payload7;
input 	write_writedata;
input 	last_write_data_8;
output 	src_payload8;
output 	src_data_33;
input 	write_writedata1;
input 	last_write_data_9;
output 	src_payload9;
input 	write_writedata2;
input 	last_write_data_10;
output 	src_payload10;
input 	write_writedata3;
input 	last_write_data_11;
output 	src_payload11;
input 	write_writedata4;
input 	last_write_data_12;
output 	src_payload12;
input 	write_writedata5;
input 	last_write_data_13;
output 	src_payload13;
input 	write_writedata6;
input 	last_write_data_14;
output 	src_payload14;
input 	write_writedata7;
input 	last_write_data_15;
output 	src_payload15;
input 	last_write_data_16;
output 	src_payload16;
output 	src_data_34;
input 	last_write_data_17;
output 	src_payload17;
input 	last_write_data_18;
output 	src_payload18;
input 	last_write_data_19;
output 	src_payload19;
input 	last_write_data_20;
output 	src_payload20;
input 	last_write_data_21;
output 	src_payload21;
input 	last_write_data_22;
output 	src_payload22;
input 	last_write_data_23;
output 	src_payload23;
input 	last_write_data_24;
output 	src_payload24;
output 	src_data_35;
input 	last_write_data_25;
output 	src_payload25;
input 	last_write_data_26;
output 	src_payload26;
input 	last_write_data_27;
output 	src_payload27;
input 	last_write_data_28;
output 	src_payload28;
input 	last_write_data_29;
output 	src_payload29;
input 	last_write_data_30;
output 	src_payload30;
input 	last_write_data_31;
output 	src_payload31;
input 	r_sync_rst;
output 	src0_valid;
input 	read_select;
output 	read_latency_shift_reg;
output 	src_data_51;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \onchip_sram_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_sram_s1_agent_rsp_fifo|mem[0][83]~q ;
wire \onchip_sram_s1_agent_rsp_fifo|mem[0][66]~q ;


Computer_System_Computer_System_mm_interconnect_2_rsp_demux rsp_demux(
	.read_latency_shift_reg_0(\onchip_sram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_83_0(\onchip_sram_s1_agent_rsp_fifo|mem[0][83]~q ),
	.mem_66_0(\onchip_sram_s1_agent_rsp_fifo|mem[0][66]~q ),
	.src0_valid1(src0_valid));

Computer_System_Computer_System_mm_interconnect_2_cmd_mux cmd_mux(
	.outclk_wire_0(outclk_wire_0),
	.readaddress_15(readaddress_15),
	.writeaddress_15(writeaddress_15),
	.q_b_0(q_b_0),
	.readaddress_2(readaddress_2),
	.writeaddress_2(writeaddress_2),
	.readaddress_3(readaddress_3),
	.writeaddress_3(writeaddress_3),
	.readaddress_4(readaddress_4),
	.writeaddress_4(writeaddress_4),
	.readaddress_5(readaddress_5),
	.writeaddress_5(writeaddress_5),
	.readaddress_6(readaddress_6),
	.writeaddress_6(writeaddress_6),
	.readaddress_7(readaddress_7),
	.writeaddress_7(writeaddress_7),
	.readaddress_8(readaddress_8),
	.writeaddress_8(writeaddress_8),
	.readaddress_9(readaddress_9),
	.writeaddress_9(writeaddress_9),
	.readaddress_10(readaddress_10),
	.writeaddress_10(writeaddress_10),
	.readaddress_11(readaddress_11),
	.writeaddress_11(writeaddress_11),
	.readaddress_12(readaddress_12),
	.writeaddress_12(writeaddress_12),
	.readaddress_13(readaddress_13),
	.writeaddress_13(writeaddress_13),
	.readaddress_14(readaddress_14),
	.writeaddress_14(writeaddress_14),
	.writeaddress_1(writeaddress_1),
	.writeaddress_0(writeaddress_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.hold_waitrequest(hold_waitrequest),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.mem_used_1(mem_used_1),
	.fifo_empty(fifo_empty),
	.last_write_collision(last_write_collision),
	.last_write_data_0(last_write_data_0),
	.control_2(control_2),
	.control_0(control_0),
	.src_payload(src_payload),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_46),
	.src_data_47(src_data_47),
	.src_data_48(src_data_48),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.src_data_32(src_data_32),
	.last_write_data_1(last_write_data_1),
	.src_payload1(src_payload1),
	.last_write_data_2(last_write_data_2),
	.src_payload2(src_payload2),
	.last_write_data_3(last_write_data_3),
	.src_payload3(src_payload3),
	.last_write_data_4(last_write_data_4),
	.src_payload4(src_payload4),
	.last_write_data_5(last_write_data_5),
	.src_payload5(src_payload5),
	.last_write_data_6(last_write_data_6),
	.src_payload6(src_payload6),
	.last_write_data_7(last_write_data_7),
	.src_payload7(src_payload7),
	.write_writedata(write_writedata),
	.last_write_data_8(last_write_data_8),
	.src_payload8(src_payload8),
	.src_data_33(src_data_33),
	.write_writedata1(write_writedata1),
	.last_write_data_9(last_write_data_9),
	.src_payload9(src_payload9),
	.write_writedata2(write_writedata2),
	.last_write_data_10(last_write_data_10),
	.src_payload10(src_payload10),
	.write_writedata3(write_writedata3),
	.last_write_data_11(last_write_data_11),
	.src_payload11(src_payload11),
	.write_writedata4(write_writedata4),
	.last_write_data_12(last_write_data_12),
	.src_payload12(src_payload12),
	.write_writedata5(write_writedata5),
	.last_write_data_13(last_write_data_13),
	.src_payload13(src_payload13),
	.write_writedata6(write_writedata6),
	.last_write_data_14(last_write_data_14),
	.src_payload14(src_payload14),
	.write_writedata7(write_writedata7),
	.last_write_data_15(last_write_data_15),
	.src_payload15(src_payload15),
	.last_write_data_16(last_write_data_16),
	.src_payload16(src_payload16),
	.src_data_34(src_data_34),
	.last_write_data_17(last_write_data_17),
	.src_payload17(src_payload17),
	.last_write_data_18(last_write_data_18),
	.src_payload18(src_payload18),
	.last_write_data_19(last_write_data_19),
	.src_payload19(src_payload19),
	.last_write_data_20(last_write_data_20),
	.src_payload20(src_payload20),
	.last_write_data_21(last_write_data_21),
	.src_payload21(src_payload21),
	.last_write_data_22(last_write_data_22),
	.src_payload22(src_payload22),
	.last_write_data_23(last_write_data_23),
	.src_payload23(src_payload23),
	.last_write_data_24(last_write_data_24),
	.src_payload24(src_payload24),
	.src_data_35(src_data_35),
	.last_write_data_25(last_write_data_25),
	.src_payload25(src_payload25),
	.last_write_data_26(last_write_data_26),
	.src_payload26(src_payload26),
	.last_write_data_27(last_write_data_27),
	.src_payload27(src_payload27),
	.last_write_data_28(last_write_data_28),
	.src_payload28(src_payload28),
	.last_write_data_29(last_write_data_29),
	.src_payload29(src_payload29),
	.last_write_data_30(last_write_data_30),
	.src_payload30(src_payload30),
	.last_write_data_31(last_write_data_31),
	.src_payload31(src_payload31),
	.r_sync_rst(r_sync_rst),
	.read_select(read_select),
	.src_data_51(src_data_51));

Computer_System_altera_avalon_sc_fifo_6 onchip_sram_s1_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.mem_used_1(mem_used_1),
	.fifo_empty(fifo_empty),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\onchip_sram_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_83_0(\onchip_sram_s1_agent_rsp_fifo|mem[0][83]~q ),
	.mem_66_0(\onchip_sram_s1_agent_rsp_fifo|mem[0][66]~q ),
	.read_select(read_select),
	.read_latency_shift_reg(read_latency_shift_reg));

Computer_System_altera_merlin_master_agent_2 dma_1_write_master_agent(
	.clk(outclk_wire_0),
	.hold_waitrequest1(hold_waitrequest),
	.r_sync_rst(r_sync_rst));

Computer_System_altera_merlin_slave_translator_2 onchip_sram_s1_translator(
	.clk(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.saved_grant_0(saved_grant_0),
	.mem_used_1(mem_used_1),
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\onchip_sram_s1_translator|read_latency_shift_reg[0]~q ),
	.read_select(read_select),
	.read_latency_shift_reg(read_latency_shift_reg));

endmodule

module Computer_System_altera_avalon_sc_fifo_6 (
	clk,
	hold_waitrequest,
	saved_grant_0,
	saved_grant_1,
	mem_used_1,
	fifo_empty,
	reset,
	read_latency_shift_reg_0,
	mem_83_0,
	mem_66_0,
	read_select,
	read_latency_shift_reg)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	hold_waitrequest;
input 	saved_grant_0;
input 	saved_grant_1;
output 	mem_used_1;
input 	fifo_empty;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_83_0;
output 	mem_66_0;
input 	read_select;
input 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][83]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][66]~q ;
wire \mem~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][83] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_83_0),
	.prn(vcc));
defparam \mem[0][83] .is_wysiwyg = "true";
defparam \mem[0][83] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!read_latency_shift_reg),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'h0FDF0FDF0FDF0FDF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!read_latency_shift_reg_0),
	.datae(!read_select),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h0F0F0F0F0F001F00;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][83] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][83]~q ),
	.prn(vcc));
defparam \mem[1][83] .is_wysiwyg = "true";
defparam \mem[1][83] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!\mem[1][83]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!saved_grant_1),
	.datab(!mem_used_1),
	.datac(!fifo_empty),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h0437043704370437;
defparam \mem~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_master_agent_2 (
	clk,
	hold_waitrequest1,
	r_sync_rst)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	hold_waitrequest1;
input 	r_sync_rst;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas hold_waitrequest(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hold_waitrequest1),
	.prn(vcc));
defparam hold_waitrequest.is_wysiwyg = "true";
defparam hold_waitrequest.power_up = "low";

endmodule

module Computer_System_altera_merlin_slave_translator_2 (
	clk,
	hold_waitrequest,
	saved_grant_0,
	mem_used_1,
	reset,
	read_latency_shift_reg_0,
	read_select,
	read_latency_shift_reg)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	hold_waitrequest;
input 	saved_grant_0;
input 	mem_used_1;
input 	reset;
output 	read_latency_shift_reg_0;
input 	read_select;
output 	read_latency_shift_reg;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!read_select),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0010001000100010;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_2_cmd_mux (
	outclk_wire_0,
	readaddress_15,
	writeaddress_15,
	q_b_0,
	readaddress_2,
	writeaddress_2,
	readaddress_3,
	writeaddress_3,
	readaddress_4,
	writeaddress_4,
	readaddress_5,
	writeaddress_5,
	readaddress_6,
	writeaddress_6,
	readaddress_7,
	writeaddress_7,
	readaddress_8,
	writeaddress_8,
	readaddress_9,
	writeaddress_9,
	readaddress_10,
	writeaddress_10,
	readaddress_11,
	writeaddress_11,
	readaddress_12,
	writeaddress_12,
	readaddress_13,
	writeaddress_13,
	readaddress_14,
	writeaddress_14,
	writeaddress_1,
	writeaddress_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	hold_waitrequest,
	saved_grant_0,
	saved_grant_1,
	mem_used_1,
	fifo_empty,
	last_write_collision,
	last_write_data_0,
	control_2,
	control_0,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	last_write_data_1,
	src_payload1,
	last_write_data_2,
	src_payload2,
	last_write_data_3,
	src_payload3,
	last_write_data_4,
	src_payload4,
	last_write_data_5,
	src_payload5,
	last_write_data_6,
	src_payload6,
	last_write_data_7,
	src_payload7,
	write_writedata,
	last_write_data_8,
	src_payload8,
	src_data_33,
	write_writedata1,
	last_write_data_9,
	src_payload9,
	write_writedata2,
	last_write_data_10,
	src_payload10,
	write_writedata3,
	last_write_data_11,
	src_payload11,
	write_writedata4,
	last_write_data_12,
	src_payload12,
	write_writedata5,
	last_write_data_13,
	src_payload13,
	write_writedata6,
	last_write_data_14,
	src_payload14,
	write_writedata7,
	last_write_data_15,
	src_payload15,
	last_write_data_16,
	src_payload16,
	src_data_34,
	last_write_data_17,
	src_payload17,
	last_write_data_18,
	src_payload18,
	last_write_data_19,
	src_payload19,
	last_write_data_20,
	src_payload20,
	last_write_data_21,
	src_payload21,
	last_write_data_22,
	src_payload22,
	last_write_data_23,
	src_payload23,
	last_write_data_24,
	src_payload24,
	src_data_35,
	last_write_data_25,
	src_payload25,
	last_write_data_26,
	src_payload26,
	last_write_data_27,
	src_payload27,
	last_write_data_28,
	src_payload28,
	last_write_data_29,
	src_payload29,
	last_write_data_30,
	src_payload30,
	last_write_data_31,
	src_payload31,
	r_sync_rst,
	read_select,
	src_data_51)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	readaddress_15;
input 	writeaddress_15;
input 	q_b_0;
input 	readaddress_2;
input 	writeaddress_2;
input 	readaddress_3;
input 	writeaddress_3;
input 	readaddress_4;
input 	writeaddress_4;
input 	readaddress_5;
input 	writeaddress_5;
input 	readaddress_6;
input 	writeaddress_6;
input 	readaddress_7;
input 	writeaddress_7;
input 	readaddress_8;
input 	writeaddress_8;
input 	readaddress_9;
input 	writeaddress_9;
input 	readaddress_10;
input 	writeaddress_10;
input 	readaddress_11;
input 	writeaddress_11;
input 	readaddress_12;
input 	writeaddress_12;
input 	readaddress_13;
input 	writeaddress_13;
input 	readaddress_14;
input 	writeaddress_14;
input 	writeaddress_1;
input 	writeaddress_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	hold_waitrequest;
output 	saved_grant_0;
output 	saved_grant_1;
input 	mem_used_1;
input 	fifo_empty;
input 	last_write_collision;
input 	last_write_data_0;
input 	control_2;
input 	control_0;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
output 	src_data_32;
input 	last_write_data_1;
output 	src_payload1;
input 	last_write_data_2;
output 	src_payload2;
input 	last_write_data_3;
output 	src_payload3;
input 	last_write_data_4;
output 	src_payload4;
input 	last_write_data_5;
output 	src_payload5;
input 	last_write_data_6;
output 	src_payload6;
input 	last_write_data_7;
output 	src_payload7;
input 	write_writedata;
input 	last_write_data_8;
output 	src_payload8;
output 	src_data_33;
input 	write_writedata1;
input 	last_write_data_9;
output 	src_payload9;
input 	write_writedata2;
input 	last_write_data_10;
output 	src_payload10;
input 	write_writedata3;
input 	last_write_data_11;
output 	src_payload11;
input 	write_writedata4;
input 	last_write_data_12;
output 	src_payload12;
input 	write_writedata5;
input 	last_write_data_13;
output 	src_payload13;
input 	write_writedata6;
input 	last_write_data_14;
output 	src_payload14;
input 	write_writedata7;
input 	last_write_data_15;
output 	src_payload15;
input 	last_write_data_16;
output 	src_payload16;
output 	src_data_34;
input 	last_write_data_17;
output 	src_payload17;
input 	last_write_data_18;
output 	src_payload18;
input 	last_write_data_19;
output 	src_payload19;
input 	last_write_data_20;
output 	src_payload20;
input 	last_write_data_21;
output 	src_payload21;
input 	last_write_data_22;
output 	src_payload22;
input 	last_write_data_23;
output 	src_payload23;
input 	last_write_data_24;
output 	src_payload24;
output 	src_data_35;
input 	last_write_data_25;
output 	src_payload25;
input 	last_write_data_26;
output 	src_payload26;
input 	last_write_data_27;
output 	src_payload27;
input 	last_write_data_28;
output 	src_payload28;
input 	last_write_data_29;
output 	src_payload29;
input 	last_write_data_30;
output 	src_payload30;
input 	last_write_data_31;
output 	src_payload31;
input 	r_sync_rst;
input 	read_select;
output 	src_data_51;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \WideOr1~0_combout ;
wire \update_grant~0_combout ;
wire \src_payload~0_combout ;


Computer_System_altera_merlin_arbitrator_8 arb(
	.clk(outclk_wire_0),
	.hold_waitrequest(hold_waitrequest),
	.fifo_empty(fifo_empty),
	.reset(r_sync_rst),
	.read_select(read_select),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~0_combout ),
	.grant_1(\arb|grant[1]~1_combout ));

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!last_write_collision),
	.datab(!last_write_data_0),
	.datac(!q_b_0),
	.datad(!\src_payload~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h001B001B001B001B;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_2),
	.datad(!writeaddress_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h0537053705370537;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_3),
	.datad(!writeaddress_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h0537053705370537;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_4),
	.datad(!writeaddress_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h0537053705370537;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_5),
	.datad(!writeaddress_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h0537053705370537;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_6),
	.datad(!writeaddress_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h0537053705370537;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_7),
	.datad(!writeaddress_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h0537053705370537;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_8),
	.datad(!writeaddress_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h0537053705370537;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_9),
	.datad(!writeaddress_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h0537053705370537;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_10),
	.datad(!writeaddress_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h0537053705370537;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_11),
	.datad(!writeaddress_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h0537053705370537;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_12),
	.datad(!writeaddress_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h0537053705370537;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_13),
	.datad(!writeaddress_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h0537053705370537;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!readaddress_14),
	.datad(!writeaddress_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h0537053705370537;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32]~0 (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32]~0 .extended_lut = "off";
defparam \src_data[32]~0 .lut_mask = 64'h7577757575757575;
defparam \src_data[32]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_1),
	.datad(!q_b_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h0123012301230123;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_2),
	.datad(!q_b_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h0123012301230123;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_3),
	.datad(!q_b_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h0123012301230123;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_4),
	.datad(!q_b_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h0123012301230123;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_5),
	.datad(!q_b_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h0123012301230123;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_6),
	.datad(!q_b_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h0123012301230123;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!last_write_collision),
	.datab(!\src_payload~0_combout ),
	.datac(!last_write_data_7),
	.datad(!q_b_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h0123012301230123;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata),
	.datae(!last_write_data_8),
	.dataf(!q_b_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h0055105540555055;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33]~1 (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33]~1 .extended_lut = "off";
defparam \src_data[33]~1 .lut_mask = 64'h7575757575777575;
defparam \src_data[33]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata1),
	.datae(!last_write_data_9),
	.dataf(!q_b_9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h0055105540555055;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata2),
	.datae(!last_write_data_10),
	.dataf(!q_b_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h0055105540555055;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata3),
	.datae(!last_write_data_11),
	.dataf(!q_b_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h0055105540555055;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata4),
	.datae(!last_write_data_12),
	.dataf(!q_b_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h0055105540555055;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata5),
	.datae(!last_write_data_13),
	.dataf(!q_b_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h0055105540555055;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata6),
	.datae(!last_write_data_14),
	.dataf(!q_b_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h0055105540555055;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata7),
	.datae(!last_write_data_15),
	.dataf(!q_b_15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h0055105540555055;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata),
	.datae(!last_write_data_16),
	.dataf(!q_b_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h0055105540555055;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34]~2 (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34]~2 .extended_lut = "off";
defparam \src_data[34]~2 .lut_mask = 64'h7575757775757575;
defparam \src_data[34]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata1),
	.datae(!last_write_data_17),
	.dataf(!q_b_17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h0055105540555055;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata2),
	.datae(!last_write_data_18),
	.dataf(!q_b_18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h0055105540555055;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata3),
	.datae(!last_write_data_19),
	.dataf(!q_b_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h0055105540555055;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata4),
	.datae(!last_write_data_20),
	.dataf(!q_b_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h0055105540555055;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata5),
	.datae(!last_write_data_21),
	.dataf(!q_b_21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h0055105540555055;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata6),
	.datae(!last_write_data_22),
	.dataf(!q_b_22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h0055105540555055;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata7),
	.datae(!last_write_data_23),
	.dataf(!q_b_23),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h0055105540555055;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata),
	.datae(!last_write_data_24),
	.dataf(!q_b_24),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h0055105540555055;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35]~3 (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!control_2),
	.datad(!control_0),
	.datae(!writeaddress_1),
	.dataf(!writeaddress_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35]~3 .extended_lut = "off";
defparam \src_data[35]~3 .lut_mask = 64'h7575757575757577;
defparam \src_data[35]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata1),
	.datae(!last_write_data_25),
	.dataf(!q_b_25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h0055105540555055;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata2),
	.datae(!last_write_data_26),
	.dataf(!q_b_26),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h0055105540555055;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata3),
	.datae(!last_write_data_27),
	.dataf(!q_b_27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h0055105540555055;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata4),
	.datae(!last_write_data_28),
	.dataf(!q_b_28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h0055105540555055;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata5),
	.datae(!last_write_data_29),
	.dataf(!q_b_29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h0055105540555055;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata6),
	.datae(!last_write_data_30),
	.dataf(!q_b_30),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h0055105540555055;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!saved_grant_1),
	.datab(!last_write_collision),
	.datac(!control_2),
	.datad(!write_writedata7),
	.datae(!last_write_data_31),
	.dataf(!q_b_31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h0055105540555055;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[51] (
	.dataa(!saved_grant_0),
	.datab(!readaddress_15),
	.datac(!saved_grant_1),
	.datad(!writeaddress_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[51] .extended_lut = "off";
defparam \src_data[51] .lut_mask = 64'h111F111F111F111F;
defparam \src_data[51] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!fifo_empty),
	.datad(!read_select),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'h0357035703570357;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!mem_used_1),
	.datae(!\packet_in_progress~q ),
	.dataf(!\WideOr1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF0000BFAA1500;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_1),
	.datab(!control_2),
	.datac(!control_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h4545454545454545;
defparam \src_payload~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_arbitrator_8 (
	clk,
	hold_waitrequest,
	fifo_empty,
	reset,
	read_select,
	grant_0,
	update_grant,
	grant_1)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	hold_waitrequest;
input 	fifo_empty;
input 	reset;
input 	read_select;
output 	grant_0;
input 	update_grant;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!hold_waitrequest),
	.datab(!fifo_empty),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!read_select),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'h0000505400005054;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!hold_waitrequest),
	.datab(!fifo_empty),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!read_select),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'h1011001110110011;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!hold_waitrequest),
	.datab(!fifo_empty),
	.datac(!read_select),
	.datad(!update_grant),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h0015001500150015;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_2_rsp_demux (
	read_latency_shift_reg_0,
	mem_83_0,
	mem_66_0,
	src0_valid1)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
input 	mem_83_0;
input 	mem_66_0;
output 	src0_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_83_0),
	.datac(!mem_66_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h5151515151515151;
defparam src0_valid.shared_arith = "off";

endmodule

module Computer_System_Computer_System_Onchip_SRAM (
	ram_block1a32,
	ram_block1a0,
	ram_block1a33,
	ram_block1a1,
	ram_block1a34,
	ram_block1a2,
	ram_block1a35,
	ram_block1a3,
	ram_block1a36,
	ram_block1a4,
	ram_block1a37,
	ram_block1a5,
	ram_block1a38,
	ram_block1a6,
	ram_block1a39,
	ram_block1a7,
	ram_block1a40,
	ram_block1a8,
	ram_block1a41,
	ram_block1a9,
	ram_block1a42,
	ram_block1a10,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a59,
	ram_block1a27,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	outclk_wire_0,
	readaddress_15,
	writeaddress_15,
	l1_w0_n0_mux_dataout,
	l1_w1_n0_mux_dataout,
	l1_w2_n0_mux_dataout,
	l1_w3_n0_mux_dataout,
	l1_w4_n0_mux_dataout,
	l1_w5_n0_mux_dataout,
	l1_w6_n0_mux_dataout,
	l1_w7_n0_mux_dataout,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w16_n0_mux_dataout,
	l1_w17_n0_mux_dataout,
	l1_w18_n0_mux_dataout,
	l1_w19_n0_mux_dataout,
	l1_w20_n0_mux_dataout,
	l1_w21_n0_mux_dataout,
	l1_w22_n0_mux_dataout,
	l1_w23_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout,
	hold_waitrequest,
	saved_grant_0,
	saved_grant_1,
	mem_used_1,
	fifo_empty,
	wren,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_data_33,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_34,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_data_35,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	address_reg_a_0,
	l1_w16_n0_mux_dataout1,
	l1_w17_n0_mux_dataout1,
	l1_w18_n0_mux_dataout1,
	l1_w19_n0_mux_dataout1,
	l1_w20_n0_mux_dataout1,
	l1_w21_n0_mux_dataout1,
	l1_w22_n0_mux_dataout1,
	l1_w23_n0_mux_dataout1,
	l1_w8_n0_mux_dataout1,
	l1_w9_n0_mux_dataout1,
	l1_w10_n0_mux_dataout1,
	l1_w11_n0_mux_dataout1,
	l1_w12_n0_mux_dataout1,
	l1_w13_n0_mux_dataout1,
	l1_w14_n0_mux_dataout1,
	l1_w15_n0_mux_dataout1,
	l1_w24_n0_mux_dataout1,
	l1_w25_n0_mux_dataout1,
	l1_w26_n0_mux_dataout1,
	l1_w27_n0_mux_dataout1,
	l1_w28_n0_mux_dataout1,
	l1_w29_n0_mux_dataout1,
	l1_w30_n0_mux_dataout1,
	l1_w31_n0_mux_dataout1,
	src_data_51,
	onchip_sram_s2_address_13,
	onchip_sram_s2_chipselect,
	onchip_sram_s2_write,
	onchip_sram_clk2_clk,
	onchip_sram_reset2_reset_req,
	onchip_sram_s2_clken,
	onchip_sram_s2_writedata_0,
	onchip_sram_s2_address_0,
	onchip_sram_s2_address_1,
	onchip_sram_s2_address_2,
	onchip_sram_s2_address_3,
	onchip_sram_s2_address_4,
	onchip_sram_s2_address_5,
	onchip_sram_s2_address_6,
	onchip_sram_s2_address_7,
	onchip_sram_s2_address_8,
	onchip_sram_s2_address_9,
	onchip_sram_s2_address_10,
	onchip_sram_s2_address_11,
	onchip_sram_s2_address_12,
	onchip_sram_s2_byteenable_0,
	onchip_sram_s2_writedata_1,
	onchip_sram_s2_writedata_2,
	onchip_sram_s2_writedata_3,
	onchip_sram_s2_writedata_4,
	onchip_sram_s2_writedata_5,
	onchip_sram_s2_writedata_6,
	onchip_sram_s2_writedata_7,
	onchip_sram_s2_writedata_8,
	onchip_sram_s2_byteenable_1,
	onchip_sram_s2_writedata_9,
	onchip_sram_s2_writedata_10,
	onchip_sram_s2_writedata_11,
	onchip_sram_s2_writedata_12,
	onchip_sram_s2_writedata_13,
	onchip_sram_s2_writedata_14,
	onchip_sram_s2_writedata_15,
	onchip_sram_s2_writedata_16,
	onchip_sram_s2_byteenable_2,
	onchip_sram_s2_writedata_17,
	onchip_sram_s2_writedata_18,
	onchip_sram_s2_writedata_19,
	onchip_sram_s2_writedata_20,
	onchip_sram_s2_writedata_21,
	onchip_sram_s2_writedata_22,
	onchip_sram_s2_writedata_23,
	onchip_sram_s2_writedata_24,
	onchip_sram_s2_byteenable_3,
	onchip_sram_s2_writedata_25,
	onchip_sram_s2_writedata_26,
	onchip_sram_s2_writedata_27,
	onchip_sram_s2_writedata_28,
	onchip_sram_s2_writedata_29,
	onchip_sram_s2_writedata_30,
	onchip_sram_s2_writedata_31)/* synthesis synthesis_greybox=0 */;
output 	ram_block1a32;
output 	ram_block1a0;
output 	ram_block1a33;
output 	ram_block1a1;
output 	ram_block1a34;
output 	ram_block1a2;
output 	ram_block1a35;
output 	ram_block1a3;
output 	ram_block1a36;
output 	ram_block1a4;
output 	ram_block1a37;
output 	ram_block1a5;
output 	ram_block1a38;
output 	ram_block1a6;
output 	ram_block1a39;
output 	ram_block1a7;
output 	ram_block1a40;
output 	ram_block1a8;
output 	ram_block1a41;
output 	ram_block1a9;
output 	ram_block1a42;
output 	ram_block1a10;
output 	ram_block1a43;
output 	ram_block1a11;
output 	ram_block1a44;
output 	ram_block1a12;
output 	ram_block1a45;
output 	ram_block1a13;
output 	ram_block1a46;
output 	ram_block1a14;
output 	ram_block1a47;
output 	ram_block1a15;
output 	ram_block1a56;
output 	ram_block1a24;
output 	ram_block1a57;
output 	ram_block1a25;
output 	ram_block1a58;
output 	ram_block1a26;
output 	ram_block1a59;
output 	ram_block1a27;
output 	ram_block1a60;
output 	ram_block1a28;
output 	ram_block1a61;
output 	ram_block1a29;
output 	ram_block1a62;
output 	ram_block1a30;
output 	ram_block1a63;
output 	ram_block1a31;
input 	outclk_wire_0;
input 	readaddress_15;
input 	writeaddress_15;
output 	l1_w0_n0_mux_dataout;
output 	l1_w1_n0_mux_dataout;
output 	l1_w2_n0_mux_dataout;
output 	l1_w3_n0_mux_dataout;
output 	l1_w4_n0_mux_dataout;
output 	l1_w5_n0_mux_dataout;
output 	l1_w6_n0_mux_dataout;
output 	l1_w7_n0_mux_dataout;
output 	l1_w8_n0_mux_dataout;
output 	l1_w9_n0_mux_dataout;
output 	l1_w10_n0_mux_dataout;
output 	l1_w11_n0_mux_dataout;
output 	l1_w12_n0_mux_dataout;
output 	l1_w13_n0_mux_dataout;
output 	l1_w14_n0_mux_dataout;
output 	l1_w15_n0_mux_dataout;
output 	l1_w16_n0_mux_dataout;
output 	l1_w17_n0_mux_dataout;
output 	l1_w18_n0_mux_dataout;
output 	l1_w19_n0_mux_dataout;
output 	l1_w20_n0_mux_dataout;
output 	l1_w21_n0_mux_dataout;
output 	l1_w22_n0_mux_dataout;
output 	l1_w23_n0_mux_dataout;
output 	l1_w24_n0_mux_dataout;
output 	l1_w25_n0_mux_dataout;
output 	l1_w26_n0_mux_dataout;
output 	l1_w27_n0_mux_dataout;
output 	l1_w28_n0_mux_dataout;
output 	l1_w29_n0_mux_dataout;
output 	l1_w30_n0_mux_dataout;
output 	l1_w31_n0_mux_dataout;
input 	hold_waitrequest;
input 	saved_grant_0;
input 	saved_grant_1;
input 	mem_used_1;
input 	fifo_empty;
output 	wren;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_data_33;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_data_34;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_data_35;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
output 	address_reg_a_0;
output 	l1_w16_n0_mux_dataout1;
output 	l1_w17_n0_mux_dataout1;
output 	l1_w18_n0_mux_dataout1;
output 	l1_w19_n0_mux_dataout1;
output 	l1_w20_n0_mux_dataout1;
output 	l1_w21_n0_mux_dataout1;
output 	l1_w22_n0_mux_dataout1;
output 	l1_w23_n0_mux_dataout1;
output 	l1_w8_n0_mux_dataout1;
output 	l1_w9_n0_mux_dataout1;
output 	l1_w10_n0_mux_dataout1;
output 	l1_w11_n0_mux_dataout1;
output 	l1_w12_n0_mux_dataout1;
output 	l1_w13_n0_mux_dataout1;
output 	l1_w14_n0_mux_dataout1;
output 	l1_w15_n0_mux_dataout1;
output 	l1_w24_n0_mux_dataout1;
output 	l1_w25_n0_mux_dataout1;
output 	l1_w26_n0_mux_dataout1;
output 	l1_w27_n0_mux_dataout1;
output 	l1_w28_n0_mux_dataout1;
output 	l1_w29_n0_mux_dataout1;
output 	l1_w30_n0_mux_dataout1;
output 	l1_w31_n0_mux_dataout1;
input 	src_data_51;
input 	onchip_sram_s2_address_13;
input 	onchip_sram_s2_chipselect;
input 	onchip_sram_s2_write;
input 	onchip_sram_clk2_clk;
input 	onchip_sram_reset2_reset_req;
input 	onchip_sram_s2_clken;
input 	onchip_sram_s2_writedata_0;
input 	onchip_sram_s2_address_0;
input 	onchip_sram_s2_address_1;
input 	onchip_sram_s2_address_2;
input 	onchip_sram_s2_address_3;
input 	onchip_sram_s2_address_4;
input 	onchip_sram_s2_address_5;
input 	onchip_sram_s2_address_6;
input 	onchip_sram_s2_address_7;
input 	onchip_sram_s2_address_8;
input 	onchip_sram_s2_address_9;
input 	onchip_sram_s2_address_10;
input 	onchip_sram_s2_address_11;
input 	onchip_sram_s2_address_12;
input 	onchip_sram_s2_byteenable_0;
input 	onchip_sram_s2_writedata_1;
input 	onchip_sram_s2_writedata_2;
input 	onchip_sram_s2_writedata_3;
input 	onchip_sram_s2_writedata_4;
input 	onchip_sram_s2_writedata_5;
input 	onchip_sram_s2_writedata_6;
input 	onchip_sram_s2_writedata_7;
input 	onchip_sram_s2_writedata_8;
input 	onchip_sram_s2_byteenable_1;
input 	onchip_sram_s2_writedata_9;
input 	onchip_sram_s2_writedata_10;
input 	onchip_sram_s2_writedata_11;
input 	onchip_sram_s2_writedata_12;
input 	onchip_sram_s2_writedata_13;
input 	onchip_sram_s2_writedata_14;
input 	onchip_sram_s2_writedata_15;
input 	onchip_sram_s2_writedata_16;
input 	onchip_sram_s2_byteenable_2;
input 	onchip_sram_s2_writedata_17;
input 	onchip_sram_s2_writedata_18;
input 	onchip_sram_s2_writedata_19;
input 	onchip_sram_s2_writedata_20;
input 	onchip_sram_s2_writedata_21;
input 	onchip_sram_s2_writedata_22;
input 	onchip_sram_s2_writedata_23;
input 	onchip_sram_s2_writedata_24;
input 	onchip_sram_s2_byteenable_3;
input 	onchip_sram_s2_writedata_25;
input 	onchip_sram_s2_writedata_26;
input 	onchip_sram_s2_writedata_27;
input 	onchip_sram_s2_writedata_28;
input 	onchip_sram_s2_writedata_29;
input 	onchip_sram_s2_writedata_30;
input 	onchip_sram_s2_writedata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clocken1~combout ;


Computer_System_altsyncram_3 the_altsyncram(
	.ram_block1a32(ram_block1a32),
	.ram_block1a0(ram_block1a0),
	.ram_block1a33(ram_block1a33),
	.ram_block1a1(ram_block1a1),
	.ram_block1a34(ram_block1a34),
	.ram_block1a2(ram_block1a2),
	.ram_block1a35(ram_block1a35),
	.ram_block1a3(ram_block1a3),
	.ram_block1a36(ram_block1a36),
	.ram_block1a4(ram_block1a4),
	.ram_block1a37(ram_block1a37),
	.ram_block1a5(ram_block1a5),
	.ram_block1a38(ram_block1a38),
	.ram_block1a6(ram_block1a6),
	.ram_block1a39(ram_block1a39),
	.ram_block1a7(ram_block1a7),
	.ram_block1a40(ram_block1a40),
	.ram_block1a8(ram_block1a8),
	.ram_block1a41(ram_block1a41),
	.ram_block1a9(ram_block1a9),
	.ram_block1a42(ram_block1a42),
	.ram_block1a10(ram_block1a10),
	.ram_block1a43(ram_block1a43),
	.ram_block1a11(ram_block1a11),
	.ram_block1a44(ram_block1a44),
	.ram_block1a12(ram_block1a12),
	.ram_block1a45(ram_block1a45),
	.ram_block1a13(ram_block1a13),
	.ram_block1a46(ram_block1a46),
	.ram_block1a14(ram_block1a14),
	.ram_block1a47(ram_block1a47),
	.ram_block1a15(ram_block1a15),
	.ram_block1a56(ram_block1a56),
	.ram_block1a24(ram_block1a24),
	.ram_block1a57(ram_block1a57),
	.ram_block1a25(ram_block1a25),
	.ram_block1a58(ram_block1a58),
	.ram_block1a26(ram_block1a26),
	.ram_block1a59(ram_block1a59),
	.ram_block1a27(ram_block1a27),
	.ram_block1a60(ram_block1a60),
	.ram_block1a28(ram_block1a28),
	.ram_block1a61(ram_block1a61),
	.ram_block1a29(ram_block1a29),
	.ram_block1a62(ram_block1a62),
	.ram_block1a30(ram_block1a30),
	.ram_block1a63(ram_block1a63),
	.ram_block1a31(ram_block1a31),
	.clock0(outclk_wire_0),
	.readaddress_15(readaddress_15),
	.writeaddress_15(writeaddress_15),
	.l1_w0_n0_mux_dataout(l1_w0_n0_mux_dataout),
	.l1_w1_n0_mux_dataout(l1_w1_n0_mux_dataout),
	.l1_w2_n0_mux_dataout(l1_w2_n0_mux_dataout),
	.l1_w3_n0_mux_dataout(l1_w3_n0_mux_dataout),
	.l1_w4_n0_mux_dataout(l1_w4_n0_mux_dataout),
	.l1_w5_n0_mux_dataout(l1_w5_n0_mux_dataout),
	.l1_w6_n0_mux_dataout(l1_w6_n0_mux_dataout),
	.l1_w7_n0_mux_dataout(l1_w7_n0_mux_dataout),
	.l1_w8_n0_mux_dataout(l1_w8_n0_mux_dataout),
	.l1_w9_n0_mux_dataout(l1_w9_n0_mux_dataout),
	.l1_w10_n0_mux_dataout(l1_w10_n0_mux_dataout),
	.l1_w11_n0_mux_dataout(l1_w11_n0_mux_dataout),
	.l1_w12_n0_mux_dataout(l1_w12_n0_mux_dataout),
	.l1_w13_n0_mux_dataout(l1_w13_n0_mux_dataout),
	.l1_w14_n0_mux_dataout(l1_w14_n0_mux_dataout),
	.l1_w15_n0_mux_dataout(l1_w15_n0_mux_dataout),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout),
	.l1_w24_n0_mux_dataout(l1_w24_n0_mux_dataout),
	.l1_w25_n0_mux_dataout(l1_w25_n0_mux_dataout),
	.l1_w26_n0_mux_dataout(l1_w26_n0_mux_dataout),
	.l1_w27_n0_mux_dataout(l1_w27_n0_mux_dataout),
	.l1_w28_n0_mux_dataout(l1_w28_n0_mux_dataout),
	.l1_w29_n0_mux_dataout(l1_w29_n0_mux_dataout),
	.l1_w30_n0_mux_dataout(l1_w30_n0_mux_dataout),
	.l1_w31_n0_mux_dataout(l1_w31_n0_mux_dataout),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.wren(wren),
	.clocken0(r_early_rst),
	.clocken1(\clocken1~combout ),
	.data_a({src_payload31,src_payload30,src_payload29,src_payload28,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,
src_payload12,src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.address_a({src_data_51,src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.address_reg_a_0(address_reg_a_0),
	.l1_w16_n0_mux_dataout1(l1_w16_n0_mux_dataout1),
	.l1_w17_n0_mux_dataout1(l1_w17_n0_mux_dataout1),
	.l1_w18_n0_mux_dataout1(l1_w18_n0_mux_dataout1),
	.l1_w19_n0_mux_dataout1(l1_w19_n0_mux_dataout1),
	.l1_w20_n0_mux_dataout1(l1_w20_n0_mux_dataout1),
	.l1_w21_n0_mux_dataout1(l1_w21_n0_mux_dataout1),
	.l1_w22_n0_mux_dataout1(l1_w22_n0_mux_dataout1),
	.l1_w23_n0_mux_dataout1(l1_w23_n0_mux_dataout1),
	.l1_w8_n0_mux_dataout1(l1_w8_n0_mux_dataout1),
	.l1_w9_n0_mux_dataout1(l1_w9_n0_mux_dataout1),
	.l1_w10_n0_mux_dataout1(l1_w10_n0_mux_dataout1),
	.l1_w11_n0_mux_dataout1(l1_w11_n0_mux_dataout1),
	.l1_w12_n0_mux_dataout1(l1_w12_n0_mux_dataout1),
	.l1_w13_n0_mux_dataout1(l1_w13_n0_mux_dataout1),
	.l1_w14_n0_mux_dataout1(l1_w14_n0_mux_dataout1),
	.l1_w15_n0_mux_dataout1(l1_w15_n0_mux_dataout1),
	.l1_w24_n0_mux_dataout1(l1_w24_n0_mux_dataout1),
	.l1_w25_n0_mux_dataout1(l1_w25_n0_mux_dataout1),
	.l1_w26_n0_mux_dataout1(l1_w26_n0_mux_dataout1),
	.l1_w27_n0_mux_dataout1(l1_w27_n0_mux_dataout1),
	.l1_w28_n0_mux_dataout1(l1_w28_n0_mux_dataout1),
	.l1_w29_n0_mux_dataout1(l1_w29_n0_mux_dataout1),
	.l1_w30_n0_mux_dataout1(l1_w30_n0_mux_dataout1),
	.l1_w31_n0_mux_dataout1(l1_w31_n0_mux_dataout1),
	.address_b({onchip_sram_s2_address_13,onchip_sram_s2_address_12,onchip_sram_s2_address_11,onchip_sram_s2_address_10,onchip_sram_s2_address_9,onchip_sram_s2_address_8,onchip_sram_s2_address_7,onchip_sram_s2_address_6,onchip_sram_s2_address_5,onchip_sram_s2_address_4,
onchip_sram_s2_address_3,onchip_sram_s2_address_2,onchip_sram_s2_address_1,onchip_sram_s2_address_0}),
	.onchip_sram_s2_chipselect(onchip_sram_s2_chipselect),
	.onchip_sram_s2_write(onchip_sram_s2_write),
	.clock1(onchip_sram_clk2_clk),
	.data_b({onchip_sram_s2_writedata_31,onchip_sram_s2_writedata_30,onchip_sram_s2_writedata_29,onchip_sram_s2_writedata_28,onchip_sram_s2_writedata_27,onchip_sram_s2_writedata_26,onchip_sram_s2_writedata_25,onchip_sram_s2_writedata_24,onchip_sram_s2_writedata_23,
onchip_sram_s2_writedata_22,onchip_sram_s2_writedata_21,onchip_sram_s2_writedata_20,onchip_sram_s2_writedata_19,onchip_sram_s2_writedata_18,onchip_sram_s2_writedata_17,onchip_sram_s2_writedata_16,onchip_sram_s2_writedata_15,onchip_sram_s2_writedata_14,
onchip_sram_s2_writedata_13,onchip_sram_s2_writedata_12,onchip_sram_s2_writedata_11,onchip_sram_s2_writedata_10,onchip_sram_s2_writedata_9,onchip_sram_s2_writedata_8,onchip_sram_s2_writedata_7,onchip_sram_s2_writedata_6,onchip_sram_s2_writedata_5,
onchip_sram_s2_writedata_4,onchip_sram_s2_writedata_3,onchip_sram_s2_writedata_2,onchip_sram_s2_writedata_1,onchip_sram_s2_writedata_0}),
	.byteena_b({onchip_sram_s2_byteenable_3,onchip_sram_s2_byteenable_2,onchip_sram_s2_byteenable_1,onchip_sram_s2_byteenable_0}));

cyclonev_lcell_comb clocken1(
	.dataa(!onchip_sram_reset2_reset_req),
	.datab(!onchip_sram_s2_clken),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clocken1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam clocken1.extended_lut = "off";
defparam clocken1.lut_mask = 64'h2222222222222222;
defparam clocken1.shared_arith = "off";

cyclonev_lcell_comb \wren~0 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_1),
	.datac(!mem_used_1),
	.datad(!fifo_empty),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wren),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'h0010001000100010;
defparam \wren~0 .shared_arith = "off";

endmodule

module Computer_System_altsyncram_3 (
	ram_block1a32,
	ram_block1a0,
	ram_block1a33,
	ram_block1a1,
	ram_block1a34,
	ram_block1a2,
	ram_block1a35,
	ram_block1a3,
	ram_block1a36,
	ram_block1a4,
	ram_block1a37,
	ram_block1a5,
	ram_block1a38,
	ram_block1a6,
	ram_block1a39,
	ram_block1a7,
	ram_block1a40,
	ram_block1a8,
	ram_block1a41,
	ram_block1a9,
	ram_block1a42,
	ram_block1a10,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a59,
	ram_block1a27,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	clock0,
	readaddress_15,
	writeaddress_15,
	l1_w0_n0_mux_dataout,
	l1_w1_n0_mux_dataout,
	l1_w2_n0_mux_dataout,
	l1_w3_n0_mux_dataout,
	l1_w4_n0_mux_dataout,
	l1_w5_n0_mux_dataout,
	l1_w6_n0_mux_dataout,
	l1_w7_n0_mux_dataout,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w16_n0_mux_dataout,
	l1_w17_n0_mux_dataout,
	l1_w18_n0_mux_dataout,
	l1_w19_n0_mux_dataout,
	l1_w20_n0_mux_dataout,
	l1_w21_n0_mux_dataout,
	l1_w22_n0_mux_dataout,
	l1_w23_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout,
	saved_grant_0,
	saved_grant_1,
	wren,
	clocken0,
	clocken1,
	data_a,
	address_a,
	byteena_a,
	address_reg_a_0,
	l1_w16_n0_mux_dataout1,
	l1_w17_n0_mux_dataout1,
	l1_w18_n0_mux_dataout1,
	l1_w19_n0_mux_dataout1,
	l1_w20_n0_mux_dataout1,
	l1_w21_n0_mux_dataout1,
	l1_w22_n0_mux_dataout1,
	l1_w23_n0_mux_dataout1,
	l1_w8_n0_mux_dataout1,
	l1_w9_n0_mux_dataout1,
	l1_w10_n0_mux_dataout1,
	l1_w11_n0_mux_dataout1,
	l1_w12_n0_mux_dataout1,
	l1_w13_n0_mux_dataout1,
	l1_w14_n0_mux_dataout1,
	l1_w15_n0_mux_dataout1,
	l1_w24_n0_mux_dataout1,
	l1_w25_n0_mux_dataout1,
	l1_w26_n0_mux_dataout1,
	l1_w27_n0_mux_dataout1,
	l1_w28_n0_mux_dataout1,
	l1_w29_n0_mux_dataout1,
	l1_w30_n0_mux_dataout1,
	l1_w31_n0_mux_dataout1,
	address_b,
	onchip_sram_s2_chipselect,
	onchip_sram_s2_write,
	clock1,
	data_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
output 	ram_block1a32;
output 	ram_block1a0;
output 	ram_block1a33;
output 	ram_block1a1;
output 	ram_block1a34;
output 	ram_block1a2;
output 	ram_block1a35;
output 	ram_block1a3;
output 	ram_block1a36;
output 	ram_block1a4;
output 	ram_block1a37;
output 	ram_block1a5;
output 	ram_block1a38;
output 	ram_block1a6;
output 	ram_block1a39;
output 	ram_block1a7;
output 	ram_block1a40;
output 	ram_block1a8;
output 	ram_block1a41;
output 	ram_block1a9;
output 	ram_block1a42;
output 	ram_block1a10;
output 	ram_block1a43;
output 	ram_block1a11;
output 	ram_block1a44;
output 	ram_block1a12;
output 	ram_block1a45;
output 	ram_block1a13;
output 	ram_block1a46;
output 	ram_block1a14;
output 	ram_block1a47;
output 	ram_block1a15;
output 	ram_block1a56;
output 	ram_block1a24;
output 	ram_block1a57;
output 	ram_block1a25;
output 	ram_block1a58;
output 	ram_block1a26;
output 	ram_block1a59;
output 	ram_block1a27;
output 	ram_block1a60;
output 	ram_block1a28;
output 	ram_block1a61;
output 	ram_block1a29;
output 	ram_block1a62;
output 	ram_block1a30;
output 	ram_block1a63;
output 	ram_block1a31;
input 	clock0;
input 	readaddress_15;
input 	writeaddress_15;
output 	l1_w0_n0_mux_dataout;
output 	l1_w1_n0_mux_dataout;
output 	l1_w2_n0_mux_dataout;
output 	l1_w3_n0_mux_dataout;
output 	l1_w4_n0_mux_dataout;
output 	l1_w5_n0_mux_dataout;
output 	l1_w6_n0_mux_dataout;
output 	l1_w7_n0_mux_dataout;
output 	l1_w8_n0_mux_dataout;
output 	l1_w9_n0_mux_dataout;
output 	l1_w10_n0_mux_dataout;
output 	l1_w11_n0_mux_dataout;
output 	l1_w12_n0_mux_dataout;
output 	l1_w13_n0_mux_dataout;
output 	l1_w14_n0_mux_dataout;
output 	l1_w15_n0_mux_dataout;
output 	l1_w16_n0_mux_dataout;
output 	l1_w17_n0_mux_dataout;
output 	l1_w18_n0_mux_dataout;
output 	l1_w19_n0_mux_dataout;
output 	l1_w20_n0_mux_dataout;
output 	l1_w21_n0_mux_dataout;
output 	l1_w22_n0_mux_dataout;
output 	l1_w23_n0_mux_dataout;
output 	l1_w24_n0_mux_dataout;
output 	l1_w25_n0_mux_dataout;
output 	l1_w26_n0_mux_dataout;
output 	l1_w27_n0_mux_dataout;
output 	l1_w28_n0_mux_dataout;
output 	l1_w29_n0_mux_dataout;
output 	l1_w30_n0_mux_dataout;
output 	l1_w31_n0_mux_dataout;
input 	saved_grant_0;
input 	saved_grant_1;
input 	wren;
input 	clocken0;
input 	clocken1;
input 	[31:0] data_a;
input 	[13:0] address_a;
input 	[3:0] byteena_a;
output 	address_reg_a_0;
output 	l1_w16_n0_mux_dataout1;
output 	l1_w17_n0_mux_dataout1;
output 	l1_w18_n0_mux_dataout1;
output 	l1_w19_n0_mux_dataout1;
output 	l1_w20_n0_mux_dataout1;
output 	l1_w21_n0_mux_dataout1;
output 	l1_w22_n0_mux_dataout1;
output 	l1_w23_n0_mux_dataout1;
output 	l1_w8_n0_mux_dataout1;
output 	l1_w9_n0_mux_dataout1;
output 	l1_w10_n0_mux_dataout1;
output 	l1_w11_n0_mux_dataout1;
output 	l1_w12_n0_mux_dataout1;
output 	l1_w13_n0_mux_dataout1;
output 	l1_w14_n0_mux_dataout1;
output 	l1_w15_n0_mux_dataout1;
output 	l1_w24_n0_mux_dataout1;
output 	l1_w25_n0_mux_dataout1;
output 	l1_w26_n0_mux_dataout1;
output 	l1_w27_n0_mux_dataout1;
output 	l1_w28_n0_mux_dataout1;
output 	l1_w29_n0_mux_dataout1;
output 	l1_w30_n0_mux_dataout1;
output 	l1_w31_n0_mux_dataout1;
input 	[13:0] address_b;
input 	onchip_sram_s2_chipselect;
input 	onchip_sram_s2_write;
input 	clock1;
input 	[31:0] data_b;
input 	[3:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altsyncram_m062 auto_generated(
	.ram_block1a321(ram_block1a32),
	.ram_block1a01(ram_block1a0),
	.ram_block1a331(ram_block1a33),
	.ram_block1a110(ram_block1a1),
	.ram_block1a341(ram_block1a34),
	.ram_block1a210(ram_block1a2),
	.ram_block1a351(ram_block1a35),
	.ram_block1a310(ram_block1a3),
	.ram_block1a361(ram_block1a36),
	.ram_block1a410(ram_block1a4),
	.ram_block1a371(ram_block1a37),
	.ram_block1a510(ram_block1a5),
	.ram_block1a381(ram_block1a38),
	.ram_block1a64(ram_block1a6),
	.ram_block1a391(ram_block1a39),
	.ram_block1a71(ram_block1a7),
	.ram_block1a401(ram_block1a40),
	.ram_block1a81(ram_block1a8),
	.ram_block1a411(ram_block1a41),
	.ram_block1a91(ram_block1a9),
	.ram_block1a421(ram_block1a42),
	.ram_block1a101(ram_block1a10),
	.ram_block1a431(ram_block1a43),
	.ram_block1a111(ram_block1a11),
	.ram_block1a441(ram_block1a44),
	.ram_block1a121(ram_block1a12),
	.ram_block1a451(ram_block1a45),
	.ram_block1a131(ram_block1a13),
	.ram_block1a461(ram_block1a46),
	.ram_block1a141(ram_block1a14),
	.ram_block1a471(ram_block1a47),
	.ram_block1a151(ram_block1a15),
	.ram_block1a561(ram_block1a56),
	.ram_block1a241(ram_block1a24),
	.ram_block1a571(ram_block1a57),
	.ram_block1a251(ram_block1a25),
	.ram_block1a581(ram_block1a58),
	.ram_block1a261(ram_block1a26),
	.ram_block1a591(ram_block1a59),
	.ram_block1a271(ram_block1a27),
	.ram_block1a601(ram_block1a60),
	.ram_block1a281(ram_block1a28),
	.ram_block1a611(ram_block1a61),
	.ram_block1a291(ram_block1a29),
	.ram_block1a621(ram_block1a62),
	.ram_block1a301(ram_block1a30),
	.ram_block1a631(ram_block1a63),
	.ram_block1a311(ram_block1a31),
	.clock0(clock0),
	.readaddress_15(readaddress_15),
	.writeaddress_15(writeaddress_15),
	.l1_w0_n0_mux_dataout(l1_w0_n0_mux_dataout),
	.l1_w1_n0_mux_dataout(l1_w1_n0_mux_dataout),
	.l1_w2_n0_mux_dataout(l1_w2_n0_mux_dataout),
	.l1_w3_n0_mux_dataout(l1_w3_n0_mux_dataout),
	.l1_w4_n0_mux_dataout(l1_w4_n0_mux_dataout),
	.l1_w5_n0_mux_dataout(l1_w5_n0_mux_dataout),
	.l1_w6_n0_mux_dataout(l1_w6_n0_mux_dataout),
	.l1_w7_n0_mux_dataout(l1_w7_n0_mux_dataout),
	.l1_w8_n0_mux_dataout(l1_w8_n0_mux_dataout),
	.l1_w9_n0_mux_dataout(l1_w9_n0_mux_dataout),
	.l1_w10_n0_mux_dataout(l1_w10_n0_mux_dataout),
	.l1_w11_n0_mux_dataout(l1_w11_n0_mux_dataout),
	.l1_w12_n0_mux_dataout(l1_w12_n0_mux_dataout),
	.l1_w13_n0_mux_dataout(l1_w13_n0_mux_dataout),
	.l1_w14_n0_mux_dataout(l1_w14_n0_mux_dataout),
	.l1_w15_n0_mux_dataout(l1_w15_n0_mux_dataout),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout),
	.l1_w24_n0_mux_dataout(l1_w24_n0_mux_dataout),
	.l1_w25_n0_mux_dataout(l1_w25_n0_mux_dataout),
	.l1_w26_n0_mux_dataout(l1_w26_n0_mux_dataout),
	.l1_w27_n0_mux_dataout(l1_w27_n0_mux_dataout),
	.l1_w28_n0_mux_dataout(l1_w28_n0_mux_dataout),
	.l1_w29_n0_mux_dataout(l1_w29_n0_mux_dataout),
	.l1_w30_n0_mux_dataout(l1_w30_n0_mux_dataout),
	.l1_w31_n0_mux_dataout(l1_w31_n0_mux_dataout),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.wren(wren),
	.clocken0(clocken0),
	.clocken1(clocken1),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.address_reg_a_0(address_reg_a_0),
	.l1_w16_n0_mux_dataout1(l1_w16_n0_mux_dataout1),
	.l1_w17_n0_mux_dataout1(l1_w17_n0_mux_dataout1),
	.l1_w18_n0_mux_dataout1(l1_w18_n0_mux_dataout1),
	.l1_w19_n0_mux_dataout1(l1_w19_n0_mux_dataout1),
	.l1_w20_n0_mux_dataout1(l1_w20_n0_mux_dataout1),
	.l1_w21_n0_mux_dataout1(l1_w21_n0_mux_dataout1),
	.l1_w22_n0_mux_dataout1(l1_w22_n0_mux_dataout1),
	.l1_w23_n0_mux_dataout1(l1_w23_n0_mux_dataout1),
	.l1_w8_n0_mux_dataout1(l1_w8_n0_mux_dataout1),
	.l1_w9_n0_mux_dataout1(l1_w9_n0_mux_dataout1),
	.l1_w10_n0_mux_dataout1(l1_w10_n0_mux_dataout1),
	.l1_w11_n0_mux_dataout1(l1_w11_n0_mux_dataout1),
	.l1_w12_n0_mux_dataout1(l1_w12_n0_mux_dataout1),
	.l1_w13_n0_mux_dataout1(l1_w13_n0_mux_dataout1),
	.l1_w14_n0_mux_dataout1(l1_w14_n0_mux_dataout1),
	.l1_w15_n0_mux_dataout1(l1_w15_n0_mux_dataout1),
	.l1_w24_n0_mux_dataout1(l1_w24_n0_mux_dataout1),
	.l1_w25_n0_mux_dataout1(l1_w25_n0_mux_dataout1),
	.l1_w26_n0_mux_dataout1(l1_w26_n0_mux_dataout1),
	.l1_w27_n0_mux_dataout1(l1_w27_n0_mux_dataout1),
	.l1_w28_n0_mux_dataout1(l1_w28_n0_mux_dataout1),
	.l1_w29_n0_mux_dataout1(l1_w29_n0_mux_dataout1),
	.l1_w30_n0_mux_dataout1(l1_w30_n0_mux_dataout1),
	.l1_w31_n0_mux_dataout1(l1_w31_n0_mux_dataout1),
	.address_b({address_b[13],address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.onchip_sram_s2_chipselect(onchip_sram_s2_chipselect),
	.onchip_sram_s2_write(onchip_sram_s2_write),
	.clock1(clock1),
	.data_b({data_b[31],data_b[30],data_b[29],data_b[28],data_b[27],data_b[26],data_b[25],data_b[24],data_b[23],data_b[22],data_b[21],data_b[20],data_b[19],data_b[18],data_b[17],data_b[16],data_b[15],data_b[14],data_b[13],data_b[12],data_b[11],data_b[10],data_b[9],data_b[8],data_b[7],data_b[6],data_b[5],data_b[4],data_b[3],data_b[2],data_b[1],data_b[0]}),
	.byteena_b({byteena_b[3],byteena_b[2],byteena_b[1],byteena_b[0]}));

endmodule

module Computer_System_altsyncram_m062 (
	ram_block1a321,
	ram_block1a01,
	ram_block1a331,
	ram_block1a110,
	ram_block1a341,
	ram_block1a210,
	ram_block1a351,
	ram_block1a310,
	ram_block1a361,
	ram_block1a410,
	ram_block1a371,
	ram_block1a510,
	ram_block1a381,
	ram_block1a64,
	ram_block1a391,
	ram_block1a71,
	ram_block1a401,
	ram_block1a81,
	ram_block1a411,
	ram_block1a91,
	ram_block1a421,
	ram_block1a101,
	ram_block1a431,
	ram_block1a111,
	ram_block1a441,
	ram_block1a121,
	ram_block1a451,
	ram_block1a131,
	ram_block1a461,
	ram_block1a141,
	ram_block1a471,
	ram_block1a151,
	ram_block1a561,
	ram_block1a241,
	ram_block1a571,
	ram_block1a251,
	ram_block1a581,
	ram_block1a261,
	ram_block1a591,
	ram_block1a271,
	ram_block1a601,
	ram_block1a281,
	ram_block1a611,
	ram_block1a291,
	ram_block1a621,
	ram_block1a301,
	ram_block1a631,
	ram_block1a311,
	clock0,
	readaddress_15,
	writeaddress_15,
	l1_w0_n0_mux_dataout,
	l1_w1_n0_mux_dataout,
	l1_w2_n0_mux_dataout,
	l1_w3_n0_mux_dataout,
	l1_w4_n0_mux_dataout,
	l1_w5_n0_mux_dataout,
	l1_w6_n0_mux_dataout,
	l1_w7_n0_mux_dataout,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w16_n0_mux_dataout,
	l1_w17_n0_mux_dataout,
	l1_w18_n0_mux_dataout,
	l1_w19_n0_mux_dataout,
	l1_w20_n0_mux_dataout,
	l1_w21_n0_mux_dataout,
	l1_w22_n0_mux_dataout,
	l1_w23_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout,
	saved_grant_0,
	saved_grant_1,
	wren,
	clocken0,
	clocken1,
	data_a,
	address_a,
	byteena_a,
	address_reg_a_0,
	l1_w16_n0_mux_dataout1,
	l1_w17_n0_mux_dataout1,
	l1_w18_n0_mux_dataout1,
	l1_w19_n0_mux_dataout1,
	l1_w20_n0_mux_dataout1,
	l1_w21_n0_mux_dataout1,
	l1_w22_n0_mux_dataout1,
	l1_w23_n0_mux_dataout1,
	l1_w8_n0_mux_dataout1,
	l1_w9_n0_mux_dataout1,
	l1_w10_n0_mux_dataout1,
	l1_w11_n0_mux_dataout1,
	l1_w12_n0_mux_dataout1,
	l1_w13_n0_mux_dataout1,
	l1_w14_n0_mux_dataout1,
	l1_w15_n0_mux_dataout1,
	l1_w24_n0_mux_dataout1,
	l1_w25_n0_mux_dataout1,
	l1_w26_n0_mux_dataout1,
	l1_w27_n0_mux_dataout1,
	l1_w28_n0_mux_dataout1,
	l1_w29_n0_mux_dataout1,
	l1_w30_n0_mux_dataout1,
	l1_w31_n0_mux_dataout1,
	address_b,
	onchip_sram_s2_chipselect,
	onchip_sram_s2_write,
	clock1,
	data_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
output 	ram_block1a321;
output 	ram_block1a01;
output 	ram_block1a331;
output 	ram_block1a110;
output 	ram_block1a341;
output 	ram_block1a210;
output 	ram_block1a351;
output 	ram_block1a310;
output 	ram_block1a361;
output 	ram_block1a410;
output 	ram_block1a371;
output 	ram_block1a510;
output 	ram_block1a381;
output 	ram_block1a64;
output 	ram_block1a391;
output 	ram_block1a71;
output 	ram_block1a401;
output 	ram_block1a81;
output 	ram_block1a411;
output 	ram_block1a91;
output 	ram_block1a421;
output 	ram_block1a101;
output 	ram_block1a431;
output 	ram_block1a111;
output 	ram_block1a441;
output 	ram_block1a121;
output 	ram_block1a451;
output 	ram_block1a131;
output 	ram_block1a461;
output 	ram_block1a141;
output 	ram_block1a471;
output 	ram_block1a151;
output 	ram_block1a561;
output 	ram_block1a241;
output 	ram_block1a571;
output 	ram_block1a251;
output 	ram_block1a581;
output 	ram_block1a261;
output 	ram_block1a591;
output 	ram_block1a271;
output 	ram_block1a601;
output 	ram_block1a281;
output 	ram_block1a611;
output 	ram_block1a291;
output 	ram_block1a621;
output 	ram_block1a301;
output 	ram_block1a631;
output 	ram_block1a311;
input 	clock0;
input 	readaddress_15;
input 	writeaddress_15;
output 	l1_w0_n0_mux_dataout;
output 	l1_w1_n0_mux_dataout;
output 	l1_w2_n0_mux_dataout;
output 	l1_w3_n0_mux_dataout;
output 	l1_w4_n0_mux_dataout;
output 	l1_w5_n0_mux_dataout;
output 	l1_w6_n0_mux_dataout;
output 	l1_w7_n0_mux_dataout;
output 	l1_w8_n0_mux_dataout;
output 	l1_w9_n0_mux_dataout;
output 	l1_w10_n0_mux_dataout;
output 	l1_w11_n0_mux_dataout;
output 	l1_w12_n0_mux_dataout;
output 	l1_w13_n0_mux_dataout;
output 	l1_w14_n0_mux_dataout;
output 	l1_w15_n0_mux_dataout;
output 	l1_w16_n0_mux_dataout;
output 	l1_w17_n0_mux_dataout;
output 	l1_w18_n0_mux_dataout;
output 	l1_w19_n0_mux_dataout;
output 	l1_w20_n0_mux_dataout;
output 	l1_w21_n0_mux_dataout;
output 	l1_w22_n0_mux_dataout;
output 	l1_w23_n0_mux_dataout;
output 	l1_w24_n0_mux_dataout;
output 	l1_w25_n0_mux_dataout;
output 	l1_w26_n0_mux_dataout;
output 	l1_w27_n0_mux_dataout;
output 	l1_w28_n0_mux_dataout;
output 	l1_w29_n0_mux_dataout;
output 	l1_w30_n0_mux_dataout;
output 	l1_w31_n0_mux_dataout;
input 	saved_grant_0;
input 	saved_grant_1;
input 	wren;
input 	clocken0;
input 	clocken1;
input 	[31:0] data_a;
input 	[13:0] address_a;
input 	[3:0] byteena_a;
output 	address_reg_a_0;
output 	l1_w16_n0_mux_dataout1;
output 	l1_w17_n0_mux_dataout1;
output 	l1_w18_n0_mux_dataout1;
output 	l1_w19_n0_mux_dataout1;
output 	l1_w20_n0_mux_dataout1;
output 	l1_w21_n0_mux_dataout1;
output 	l1_w22_n0_mux_dataout1;
output 	l1_w23_n0_mux_dataout1;
output 	l1_w8_n0_mux_dataout1;
output 	l1_w9_n0_mux_dataout1;
output 	l1_w10_n0_mux_dataout1;
output 	l1_w11_n0_mux_dataout1;
output 	l1_w12_n0_mux_dataout1;
output 	l1_w13_n0_mux_dataout1;
output 	l1_w14_n0_mux_dataout1;
output 	l1_w15_n0_mux_dataout1;
output 	l1_w24_n0_mux_dataout1;
output 	l1_w25_n0_mux_dataout1;
output 	l1_w26_n0_mux_dataout1;
output 	l1_w27_n0_mux_dataout1;
output 	l1_w28_n0_mux_dataout1;
output 	l1_w29_n0_mux_dataout1;
output 	l1_w30_n0_mux_dataout1;
output 	l1_w31_n0_mux_dataout1;
input 	[13:0] address_b;
input 	onchip_sram_s2_chipselect;
input 	onchip_sram_s2_write;
input 	clock1;
input 	[31:0] data_b;
input 	[3:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_block1a48~portadataout ;
wire \ram_block1a48~PORTBDATAOUT0 ;
wire \ram_block1a16~portadataout ;
wire \ram_block1a16~PORTBDATAOUT0 ;
wire \ram_block1a49~portadataout ;
wire \ram_block1a49~PORTBDATAOUT0 ;
wire \ram_block1a17~portadataout ;
wire \ram_block1a17~PORTBDATAOUT0 ;
wire \ram_block1a50~portadataout ;
wire \ram_block1a50~PORTBDATAOUT0 ;
wire \ram_block1a18~portadataout ;
wire \ram_block1a18~PORTBDATAOUT0 ;
wire \ram_block1a51~portadataout ;
wire \ram_block1a51~PORTBDATAOUT0 ;
wire \ram_block1a19~portadataout ;
wire \ram_block1a19~PORTBDATAOUT0 ;
wire \ram_block1a52~portadataout ;
wire \ram_block1a52~PORTBDATAOUT0 ;
wire \ram_block1a20~portadataout ;
wire \ram_block1a20~PORTBDATAOUT0 ;
wire \ram_block1a53~portadataout ;
wire \ram_block1a53~PORTBDATAOUT0 ;
wire \ram_block1a21~portadataout ;
wire \ram_block1a21~PORTBDATAOUT0 ;
wire \ram_block1a54~portadataout ;
wire \ram_block1a54~PORTBDATAOUT0 ;
wire \ram_block1a22~portadataout ;
wire \ram_block1a22~PORTBDATAOUT0 ;
wire \ram_block1a55~portadataout ;
wire \ram_block1a55~PORTBDATAOUT0 ;
wire \ram_block1a23~portadataout ;
wire \ram_block1a23~PORTBDATAOUT0 ;
wire \address_reg_b[0]~q ;
wire \decode2|eq_node[1]~combout ;
wire \decode3|eq_node[1]~0_combout ;
wire \decode2|eq_node[0]~combout ;
wire \decode3|eq_node[0]~1_combout ;
wire \ram_block1a32~PORTBDATAOUT0 ;
wire \ram_block1a0~PORTBDATAOUT0 ;
wire \ram_block1a33~PORTBDATAOUT0 ;
wire \ram_block1a1~PORTBDATAOUT0 ;
wire \ram_block1a34~PORTBDATAOUT0 ;
wire \ram_block1a2~PORTBDATAOUT0 ;
wire \ram_block1a35~PORTBDATAOUT0 ;
wire \ram_block1a3~PORTBDATAOUT0 ;
wire \ram_block1a36~PORTBDATAOUT0 ;
wire \ram_block1a4~PORTBDATAOUT0 ;
wire \ram_block1a37~PORTBDATAOUT0 ;
wire \ram_block1a5~PORTBDATAOUT0 ;
wire \ram_block1a38~PORTBDATAOUT0 ;
wire \ram_block1a6~PORTBDATAOUT0 ;
wire \ram_block1a39~PORTBDATAOUT0 ;
wire \ram_block1a7~PORTBDATAOUT0 ;
wire \ram_block1a40~PORTBDATAOUT0 ;
wire \ram_block1a8~PORTBDATAOUT0 ;
wire \ram_block1a41~PORTBDATAOUT0 ;
wire \ram_block1a9~PORTBDATAOUT0 ;
wire \ram_block1a42~PORTBDATAOUT0 ;
wire \ram_block1a10~PORTBDATAOUT0 ;
wire \ram_block1a43~PORTBDATAOUT0 ;
wire \ram_block1a11~PORTBDATAOUT0 ;
wire \ram_block1a44~PORTBDATAOUT0 ;
wire \ram_block1a12~PORTBDATAOUT0 ;
wire \ram_block1a45~PORTBDATAOUT0 ;
wire \ram_block1a13~PORTBDATAOUT0 ;
wire \ram_block1a46~PORTBDATAOUT0 ;
wire \ram_block1a14~PORTBDATAOUT0 ;
wire \ram_block1a47~PORTBDATAOUT0 ;
wire \ram_block1a15~PORTBDATAOUT0 ;
wire \ram_block1a56~PORTBDATAOUT0 ;
wire \ram_block1a24~PORTBDATAOUT0 ;
wire \ram_block1a57~PORTBDATAOUT0 ;
wire \ram_block1a25~PORTBDATAOUT0 ;
wire \ram_block1a58~PORTBDATAOUT0 ;
wire \ram_block1a26~PORTBDATAOUT0 ;
wire \ram_block1a59~PORTBDATAOUT0 ;
wire \ram_block1a27~PORTBDATAOUT0 ;
wire \ram_block1a60~PORTBDATAOUT0 ;
wire \ram_block1a28~PORTBDATAOUT0 ;
wire \ram_block1a61~PORTBDATAOUT0 ;
wire \ram_block1a29~PORTBDATAOUT0 ;
wire \ram_block1a62~PORTBDATAOUT0 ;
wire \ram_block1a30~PORTBDATAOUT0 ;
wire \ram_block1a63~PORTBDATAOUT0 ;
wire \ram_block1a31~PORTBDATAOUT0 ;

wire [143:0] ram_block1a32_PORTADATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTADATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a34_PORTADATAOUT_bus;
wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTADATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTADATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTADATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a38_PORTADATAOUT_bus;
wire [143:0] ram_block1a38_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a39_PORTADATAOUT_bus;
wire [143:0] ram_block1a39_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a40_PORTADATAOUT_bus;
wire [143:0] ram_block1a40_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a41_PORTADATAOUT_bus;
wire [143:0] ram_block1a41_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a42_PORTADATAOUT_bus;
wire [143:0] ram_block1a42_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a43_PORTADATAOUT_bus;
wire [143:0] ram_block1a43_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a44_PORTADATAOUT_bus;
wire [143:0] ram_block1a44_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a45_PORTADATAOUT_bus;
wire [143:0] ram_block1a45_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a46_PORTADATAOUT_bus;
wire [143:0] ram_block1a46_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a47_PORTADATAOUT_bus;
wire [143:0] ram_block1a47_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a48_PORTADATAOUT_bus;
wire [143:0] ram_block1a48_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a49_PORTADATAOUT_bus;
wire [143:0] ram_block1a49_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a50_PORTADATAOUT_bus;
wire [143:0] ram_block1a50_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a51_PORTADATAOUT_bus;
wire [143:0] ram_block1a51_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a52_PORTADATAOUT_bus;
wire [143:0] ram_block1a52_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a53_PORTADATAOUT_bus;
wire [143:0] ram_block1a53_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a54_PORTADATAOUT_bus;
wire [143:0] ram_block1a54_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a55_PORTADATAOUT_bus;
wire [143:0] ram_block1a55_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a56_PORTADATAOUT_bus;
wire [143:0] ram_block1a56_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a57_PORTADATAOUT_bus;
wire [143:0] ram_block1a57_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a58_PORTADATAOUT_bus;
wire [143:0] ram_block1a58_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a59_PORTADATAOUT_bus;
wire [143:0] ram_block1a59_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a60_PORTADATAOUT_bus;
wire [143:0] ram_block1a60_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a61_PORTADATAOUT_bus;
wire [143:0] ram_block1a61_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a62_PORTADATAOUT_bus;
wire [143:0] ram_block1a62_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a63_PORTADATAOUT_bus;
wire [143:0] ram_block1a63_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign ram_block1a321 = ram_block1a32_PORTADATAOUT_bus[0];

assign \ram_block1a32~PORTBDATAOUT0  = ram_block1a32_PORTBDATAOUT_bus[0];

assign ram_block1a01 = ram_block1a0_PORTADATAOUT_bus[0];

assign \ram_block1a0~PORTBDATAOUT0  = ram_block1a0_PORTBDATAOUT_bus[0];

assign ram_block1a331 = ram_block1a33_PORTADATAOUT_bus[0];

assign \ram_block1a33~PORTBDATAOUT0  = ram_block1a33_PORTBDATAOUT_bus[0];

assign ram_block1a110 = ram_block1a1_PORTADATAOUT_bus[0];

assign \ram_block1a1~PORTBDATAOUT0  = ram_block1a1_PORTBDATAOUT_bus[0];

assign ram_block1a341 = ram_block1a34_PORTADATAOUT_bus[0];

assign \ram_block1a34~PORTBDATAOUT0  = ram_block1a34_PORTBDATAOUT_bus[0];

assign ram_block1a210 = ram_block1a2_PORTADATAOUT_bus[0];

assign \ram_block1a2~PORTBDATAOUT0  = ram_block1a2_PORTBDATAOUT_bus[0];

assign ram_block1a351 = ram_block1a35_PORTADATAOUT_bus[0];

assign \ram_block1a35~PORTBDATAOUT0  = ram_block1a35_PORTBDATAOUT_bus[0];

assign ram_block1a310 = ram_block1a3_PORTADATAOUT_bus[0];

assign \ram_block1a3~PORTBDATAOUT0  = ram_block1a3_PORTBDATAOUT_bus[0];

assign ram_block1a361 = ram_block1a36_PORTADATAOUT_bus[0];

assign \ram_block1a36~PORTBDATAOUT0  = ram_block1a36_PORTBDATAOUT_bus[0];

assign ram_block1a410 = ram_block1a4_PORTADATAOUT_bus[0];

assign \ram_block1a4~PORTBDATAOUT0  = ram_block1a4_PORTBDATAOUT_bus[0];

assign ram_block1a371 = ram_block1a37_PORTADATAOUT_bus[0];

assign \ram_block1a37~PORTBDATAOUT0  = ram_block1a37_PORTBDATAOUT_bus[0];

assign ram_block1a510 = ram_block1a5_PORTADATAOUT_bus[0];

assign \ram_block1a5~PORTBDATAOUT0  = ram_block1a5_PORTBDATAOUT_bus[0];

assign ram_block1a381 = ram_block1a38_PORTADATAOUT_bus[0];

assign \ram_block1a38~PORTBDATAOUT0  = ram_block1a38_PORTBDATAOUT_bus[0];

assign ram_block1a64 = ram_block1a6_PORTADATAOUT_bus[0];

assign \ram_block1a6~PORTBDATAOUT0  = ram_block1a6_PORTBDATAOUT_bus[0];

assign ram_block1a391 = ram_block1a39_PORTADATAOUT_bus[0];

assign \ram_block1a39~PORTBDATAOUT0  = ram_block1a39_PORTBDATAOUT_bus[0];

assign ram_block1a71 = ram_block1a7_PORTADATAOUT_bus[0];

assign \ram_block1a7~PORTBDATAOUT0  = ram_block1a7_PORTBDATAOUT_bus[0];

assign ram_block1a401 = ram_block1a40_PORTADATAOUT_bus[0];

assign \ram_block1a40~PORTBDATAOUT0  = ram_block1a40_PORTBDATAOUT_bus[0];

assign ram_block1a81 = ram_block1a8_PORTADATAOUT_bus[0];

assign \ram_block1a8~PORTBDATAOUT0  = ram_block1a8_PORTBDATAOUT_bus[0];

assign ram_block1a411 = ram_block1a41_PORTADATAOUT_bus[0];

assign \ram_block1a41~PORTBDATAOUT0  = ram_block1a41_PORTBDATAOUT_bus[0];

assign ram_block1a91 = ram_block1a9_PORTADATAOUT_bus[0];

assign \ram_block1a9~PORTBDATAOUT0  = ram_block1a9_PORTBDATAOUT_bus[0];

assign ram_block1a421 = ram_block1a42_PORTADATAOUT_bus[0];

assign \ram_block1a42~PORTBDATAOUT0  = ram_block1a42_PORTBDATAOUT_bus[0];

assign ram_block1a101 = ram_block1a10_PORTADATAOUT_bus[0];

assign \ram_block1a10~PORTBDATAOUT0  = ram_block1a10_PORTBDATAOUT_bus[0];

assign ram_block1a431 = ram_block1a43_PORTADATAOUT_bus[0];

assign \ram_block1a43~PORTBDATAOUT0  = ram_block1a43_PORTBDATAOUT_bus[0];

assign ram_block1a111 = ram_block1a11_PORTADATAOUT_bus[0];

assign \ram_block1a11~PORTBDATAOUT0  = ram_block1a11_PORTBDATAOUT_bus[0];

assign ram_block1a441 = ram_block1a44_PORTADATAOUT_bus[0];

assign \ram_block1a44~PORTBDATAOUT0  = ram_block1a44_PORTBDATAOUT_bus[0];

assign ram_block1a121 = ram_block1a12_PORTADATAOUT_bus[0];

assign \ram_block1a12~PORTBDATAOUT0  = ram_block1a12_PORTBDATAOUT_bus[0];

assign ram_block1a451 = ram_block1a45_PORTADATAOUT_bus[0];

assign \ram_block1a45~PORTBDATAOUT0  = ram_block1a45_PORTBDATAOUT_bus[0];

assign ram_block1a131 = ram_block1a13_PORTADATAOUT_bus[0];

assign \ram_block1a13~PORTBDATAOUT0  = ram_block1a13_PORTBDATAOUT_bus[0];

assign ram_block1a461 = ram_block1a46_PORTADATAOUT_bus[0];

assign \ram_block1a46~PORTBDATAOUT0  = ram_block1a46_PORTBDATAOUT_bus[0];

assign ram_block1a141 = ram_block1a14_PORTADATAOUT_bus[0];

assign \ram_block1a14~PORTBDATAOUT0  = ram_block1a14_PORTBDATAOUT_bus[0];

assign ram_block1a471 = ram_block1a47_PORTADATAOUT_bus[0];

assign \ram_block1a47~PORTBDATAOUT0  = ram_block1a47_PORTBDATAOUT_bus[0];

assign ram_block1a151 = ram_block1a15_PORTADATAOUT_bus[0];

assign \ram_block1a15~PORTBDATAOUT0  = ram_block1a15_PORTBDATAOUT_bus[0];

assign \ram_block1a48~portadataout  = ram_block1a48_PORTADATAOUT_bus[0];

assign \ram_block1a48~PORTBDATAOUT0  = ram_block1a48_PORTBDATAOUT_bus[0];

assign \ram_block1a16~portadataout  = ram_block1a16_PORTADATAOUT_bus[0];

assign \ram_block1a16~PORTBDATAOUT0  = ram_block1a16_PORTBDATAOUT_bus[0];

assign \ram_block1a49~portadataout  = ram_block1a49_PORTADATAOUT_bus[0];

assign \ram_block1a49~PORTBDATAOUT0  = ram_block1a49_PORTBDATAOUT_bus[0];

assign \ram_block1a17~portadataout  = ram_block1a17_PORTADATAOUT_bus[0];

assign \ram_block1a17~PORTBDATAOUT0  = ram_block1a17_PORTBDATAOUT_bus[0];

assign \ram_block1a50~portadataout  = ram_block1a50_PORTADATAOUT_bus[0];

assign \ram_block1a50~PORTBDATAOUT0  = ram_block1a50_PORTBDATAOUT_bus[0];

assign \ram_block1a18~portadataout  = ram_block1a18_PORTADATAOUT_bus[0];

assign \ram_block1a18~PORTBDATAOUT0  = ram_block1a18_PORTBDATAOUT_bus[0];

assign \ram_block1a51~portadataout  = ram_block1a51_PORTADATAOUT_bus[0];

assign \ram_block1a51~PORTBDATAOUT0  = ram_block1a51_PORTBDATAOUT_bus[0];

assign \ram_block1a19~portadataout  = ram_block1a19_PORTADATAOUT_bus[0];

assign \ram_block1a19~PORTBDATAOUT0  = ram_block1a19_PORTBDATAOUT_bus[0];

assign \ram_block1a52~portadataout  = ram_block1a52_PORTADATAOUT_bus[0];

assign \ram_block1a52~PORTBDATAOUT0  = ram_block1a52_PORTBDATAOUT_bus[0];

assign \ram_block1a20~portadataout  = ram_block1a20_PORTADATAOUT_bus[0];

assign \ram_block1a20~PORTBDATAOUT0  = ram_block1a20_PORTBDATAOUT_bus[0];

assign \ram_block1a53~portadataout  = ram_block1a53_PORTADATAOUT_bus[0];

assign \ram_block1a53~PORTBDATAOUT0  = ram_block1a53_PORTBDATAOUT_bus[0];

assign \ram_block1a21~portadataout  = ram_block1a21_PORTADATAOUT_bus[0];

assign \ram_block1a21~PORTBDATAOUT0  = ram_block1a21_PORTBDATAOUT_bus[0];

assign \ram_block1a54~portadataout  = ram_block1a54_PORTADATAOUT_bus[0];

assign \ram_block1a54~PORTBDATAOUT0  = ram_block1a54_PORTBDATAOUT_bus[0];

assign \ram_block1a22~portadataout  = ram_block1a22_PORTADATAOUT_bus[0];

assign \ram_block1a22~PORTBDATAOUT0  = ram_block1a22_PORTBDATAOUT_bus[0];

assign \ram_block1a55~portadataout  = ram_block1a55_PORTADATAOUT_bus[0];

assign \ram_block1a55~PORTBDATAOUT0  = ram_block1a55_PORTBDATAOUT_bus[0];

assign \ram_block1a23~portadataout  = ram_block1a23_PORTADATAOUT_bus[0];

assign \ram_block1a23~PORTBDATAOUT0  = ram_block1a23_PORTBDATAOUT_bus[0];

assign ram_block1a561 = ram_block1a56_PORTADATAOUT_bus[0];

assign \ram_block1a56~PORTBDATAOUT0  = ram_block1a56_PORTBDATAOUT_bus[0];

assign ram_block1a241 = ram_block1a24_PORTADATAOUT_bus[0];

assign \ram_block1a24~PORTBDATAOUT0  = ram_block1a24_PORTBDATAOUT_bus[0];

assign ram_block1a571 = ram_block1a57_PORTADATAOUT_bus[0];

assign \ram_block1a57~PORTBDATAOUT0  = ram_block1a57_PORTBDATAOUT_bus[0];

assign ram_block1a251 = ram_block1a25_PORTADATAOUT_bus[0];

assign \ram_block1a25~PORTBDATAOUT0  = ram_block1a25_PORTBDATAOUT_bus[0];

assign ram_block1a581 = ram_block1a58_PORTADATAOUT_bus[0];

assign \ram_block1a58~PORTBDATAOUT0  = ram_block1a58_PORTBDATAOUT_bus[0];

assign ram_block1a261 = ram_block1a26_PORTADATAOUT_bus[0];

assign \ram_block1a26~PORTBDATAOUT0  = ram_block1a26_PORTBDATAOUT_bus[0];

assign ram_block1a591 = ram_block1a59_PORTADATAOUT_bus[0];

assign \ram_block1a59~PORTBDATAOUT0  = ram_block1a59_PORTBDATAOUT_bus[0];

assign ram_block1a271 = ram_block1a27_PORTADATAOUT_bus[0];

assign \ram_block1a27~PORTBDATAOUT0  = ram_block1a27_PORTBDATAOUT_bus[0];

assign ram_block1a601 = ram_block1a60_PORTADATAOUT_bus[0];

assign \ram_block1a60~PORTBDATAOUT0  = ram_block1a60_PORTBDATAOUT_bus[0];

assign ram_block1a281 = ram_block1a28_PORTADATAOUT_bus[0];

assign \ram_block1a28~PORTBDATAOUT0  = ram_block1a28_PORTBDATAOUT_bus[0];

assign ram_block1a611 = ram_block1a61_PORTADATAOUT_bus[0];

assign \ram_block1a61~PORTBDATAOUT0  = ram_block1a61_PORTBDATAOUT_bus[0];

assign ram_block1a291 = ram_block1a29_PORTADATAOUT_bus[0];

assign \ram_block1a29~PORTBDATAOUT0  = ram_block1a29_PORTBDATAOUT_bus[0];

assign ram_block1a621 = ram_block1a62_PORTADATAOUT_bus[0];

assign \ram_block1a62~PORTBDATAOUT0  = ram_block1a62_PORTBDATAOUT_bus[0];

assign ram_block1a301 = ram_block1a30_PORTADATAOUT_bus[0];

assign \ram_block1a30~PORTBDATAOUT0  = ram_block1a30_PORTBDATAOUT_bus[0];

assign ram_block1a631 = ram_block1a63_PORTADATAOUT_bus[0];

assign \ram_block1a63~PORTBDATAOUT0  = ram_block1a63_PORTBDATAOUT_bus[0];

assign ram_block1a311 = ram_block1a31_PORTADATAOUT_bus[0];

assign \ram_block1a31~PORTBDATAOUT0  = ram_block1a31_PORTBDATAOUT_bus[0];

Computer_System_mux_2hb_1 mux5(
	.ram_block1a32(\ram_block1a32~PORTBDATAOUT0 ),
	.ram_block1a0(\ram_block1a0~PORTBDATAOUT0 ),
	.ram_block1a33(\ram_block1a33~PORTBDATAOUT0 ),
	.ram_block1a1(\ram_block1a1~PORTBDATAOUT0 ),
	.ram_block1a34(\ram_block1a34~PORTBDATAOUT0 ),
	.ram_block1a2(\ram_block1a2~PORTBDATAOUT0 ),
	.ram_block1a35(\ram_block1a35~PORTBDATAOUT0 ),
	.ram_block1a3(\ram_block1a3~PORTBDATAOUT0 ),
	.ram_block1a36(\ram_block1a36~PORTBDATAOUT0 ),
	.ram_block1a4(\ram_block1a4~PORTBDATAOUT0 ),
	.ram_block1a37(\ram_block1a37~PORTBDATAOUT0 ),
	.ram_block1a5(\ram_block1a5~PORTBDATAOUT0 ),
	.ram_block1a38(\ram_block1a38~PORTBDATAOUT0 ),
	.ram_block1a6(\ram_block1a6~PORTBDATAOUT0 ),
	.ram_block1a39(\ram_block1a39~PORTBDATAOUT0 ),
	.ram_block1a7(\ram_block1a7~PORTBDATAOUT0 ),
	.ram_block1a40(\ram_block1a40~PORTBDATAOUT0 ),
	.ram_block1a8(\ram_block1a8~PORTBDATAOUT0 ),
	.ram_block1a41(\ram_block1a41~PORTBDATAOUT0 ),
	.ram_block1a9(\ram_block1a9~PORTBDATAOUT0 ),
	.ram_block1a42(\ram_block1a42~PORTBDATAOUT0 ),
	.ram_block1a10(\ram_block1a10~PORTBDATAOUT0 ),
	.ram_block1a43(\ram_block1a43~PORTBDATAOUT0 ),
	.ram_block1a11(\ram_block1a11~PORTBDATAOUT0 ),
	.ram_block1a44(\ram_block1a44~PORTBDATAOUT0 ),
	.ram_block1a12(\ram_block1a12~PORTBDATAOUT0 ),
	.ram_block1a45(\ram_block1a45~PORTBDATAOUT0 ),
	.ram_block1a13(\ram_block1a13~PORTBDATAOUT0 ),
	.ram_block1a46(\ram_block1a46~PORTBDATAOUT0 ),
	.ram_block1a14(\ram_block1a14~PORTBDATAOUT0 ),
	.ram_block1a47(\ram_block1a47~PORTBDATAOUT0 ),
	.ram_block1a15(\ram_block1a15~PORTBDATAOUT0 ),
	.ram_block1a48(\ram_block1a48~PORTBDATAOUT0 ),
	.ram_block1a16(\ram_block1a16~PORTBDATAOUT0 ),
	.ram_block1a49(\ram_block1a49~PORTBDATAOUT0 ),
	.ram_block1a17(\ram_block1a17~PORTBDATAOUT0 ),
	.ram_block1a50(\ram_block1a50~PORTBDATAOUT0 ),
	.ram_block1a18(\ram_block1a18~PORTBDATAOUT0 ),
	.ram_block1a51(\ram_block1a51~PORTBDATAOUT0 ),
	.ram_block1a19(\ram_block1a19~PORTBDATAOUT0 ),
	.ram_block1a52(\ram_block1a52~PORTBDATAOUT0 ),
	.ram_block1a20(\ram_block1a20~PORTBDATAOUT0 ),
	.ram_block1a53(\ram_block1a53~PORTBDATAOUT0 ),
	.ram_block1a21(\ram_block1a21~PORTBDATAOUT0 ),
	.ram_block1a54(\ram_block1a54~PORTBDATAOUT0 ),
	.ram_block1a22(\ram_block1a22~PORTBDATAOUT0 ),
	.ram_block1a55(\ram_block1a55~PORTBDATAOUT0 ),
	.ram_block1a23(\ram_block1a23~PORTBDATAOUT0 ),
	.ram_block1a56(\ram_block1a56~PORTBDATAOUT0 ),
	.ram_block1a24(\ram_block1a24~PORTBDATAOUT0 ),
	.ram_block1a57(\ram_block1a57~PORTBDATAOUT0 ),
	.ram_block1a25(\ram_block1a25~PORTBDATAOUT0 ),
	.ram_block1a58(\ram_block1a58~PORTBDATAOUT0 ),
	.ram_block1a26(\ram_block1a26~PORTBDATAOUT0 ),
	.ram_block1a59(\ram_block1a59~PORTBDATAOUT0 ),
	.ram_block1a27(\ram_block1a27~PORTBDATAOUT0 ),
	.ram_block1a60(\ram_block1a60~PORTBDATAOUT0 ),
	.ram_block1a28(\ram_block1a28~PORTBDATAOUT0 ),
	.ram_block1a61(\ram_block1a61~PORTBDATAOUT0 ),
	.ram_block1a29(\ram_block1a29~PORTBDATAOUT0 ),
	.ram_block1a62(\ram_block1a62~PORTBDATAOUT0 ),
	.ram_block1a30(\ram_block1a30~PORTBDATAOUT0 ),
	.ram_block1a63(\ram_block1a63~PORTBDATAOUT0 ),
	.ram_block1a31(\ram_block1a31~PORTBDATAOUT0 ),
	.address_reg_b_0(\address_reg_b[0]~q ),
	.l1_w0_n0_mux_dataout(l1_w0_n0_mux_dataout),
	.l1_w1_n0_mux_dataout(l1_w1_n0_mux_dataout),
	.l1_w2_n0_mux_dataout(l1_w2_n0_mux_dataout),
	.l1_w3_n0_mux_dataout(l1_w3_n0_mux_dataout),
	.l1_w4_n0_mux_dataout(l1_w4_n0_mux_dataout),
	.l1_w5_n0_mux_dataout(l1_w5_n0_mux_dataout),
	.l1_w6_n0_mux_dataout(l1_w6_n0_mux_dataout),
	.l1_w7_n0_mux_dataout(l1_w7_n0_mux_dataout),
	.l1_w8_n0_mux_dataout(l1_w8_n0_mux_dataout),
	.l1_w9_n0_mux_dataout(l1_w9_n0_mux_dataout),
	.l1_w10_n0_mux_dataout(l1_w10_n0_mux_dataout),
	.l1_w11_n0_mux_dataout(l1_w11_n0_mux_dataout),
	.l1_w12_n0_mux_dataout(l1_w12_n0_mux_dataout),
	.l1_w13_n0_mux_dataout(l1_w13_n0_mux_dataout),
	.l1_w14_n0_mux_dataout(l1_w14_n0_mux_dataout),
	.l1_w15_n0_mux_dataout(l1_w15_n0_mux_dataout),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout),
	.l1_w24_n0_mux_dataout(l1_w24_n0_mux_dataout),
	.l1_w25_n0_mux_dataout(l1_w25_n0_mux_dataout),
	.l1_w26_n0_mux_dataout(l1_w26_n0_mux_dataout),
	.l1_w27_n0_mux_dataout(l1_w27_n0_mux_dataout),
	.l1_w28_n0_mux_dataout(l1_w28_n0_mux_dataout),
	.l1_w29_n0_mux_dataout(l1_w29_n0_mux_dataout),
	.l1_w30_n0_mux_dataout(l1_w30_n0_mux_dataout),
	.l1_w31_n0_mux_dataout(l1_w31_n0_mux_dataout));

Computer_System_mux_2hb mux4(
	.ram_block1a40(ram_block1a401),
	.ram_block1a8(ram_block1a81),
	.ram_block1a41(ram_block1a411),
	.ram_block1a9(ram_block1a91),
	.ram_block1a42(ram_block1a421),
	.ram_block1a10(ram_block1a101),
	.ram_block1a43(ram_block1a431),
	.ram_block1a11(ram_block1a111),
	.ram_block1a44(ram_block1a441),
	.ram_block1a12(ram_block1a121),
	.ram_block1a45(ram_block1a451),
	.ram_block1a13(ram_block1a131),
	.ram_block1a46(ram_block1a461),
	.ram_block1a14(ram_block1a141),
	.ram_block1a47(ram_block1a471),
	.ram_block1a15(ram_block1a151),
	.ram_block1a48(\ram_block1a48~portadataout ),
	.ram_block1a16(\ram_block1a16~portadataout ),
	.ram_block1a49(\ram_block1a49~portadataout ),
	.ram_block1a17(\ram_block1a17~portadataout ),
	.ram_block1a50(\ram_block1a50~portadataout ),
	.ram_block1a18(\ram_block1a18~portadataout ),
	.ram_block1a51(\ram_block1a51~portadataout ),
	.ram_block1a19(\ram_block1a19~portadataout ),
	.ram_block1a52(\ram_block1a52~portadataout ),
	.ram_block1a20(\ram_block1a20~portadataout ),
	.ram_block1a53(\ram_block1a53~portadataout ),
	.ram_block1a21(\ram_block1a21~portadataout ),
	.ram_block1a54(\ram_block1a54~portadataout ),
	.ram_block1a22(\ram_block1a22~portadataout ),
	.ram_block1a55(\ram_block1a55~portadataout ),
	.ram_block1a23(\ram_block1a23~portadataout ),
	.ram_block1a56(ram_block1a561),
	.ram_block1a24(ram_block1a241),
	.ram_block1a57(ram_block1a571),
	.ram_block1a25(ram_block1a251),
	.ram_block1a58(ram_block1a581),
	.ram_block1a26(ram_block1a261),
	.ram_block1a59(ram_block1a591),
	.ram_block1a27(ram_block1a271),
	.ram_block1a60(ram_block1a601),
	.ram_block1a28(ram_block1a281),
	.ram_block1a61(ram_block1a611),
	.ram_block1a29(ram_block1a291),
	.ram_block1a62(ram_block1a621),
	.ram_block1a30(ram_block1a301),
	.ram_block1a63(ram_block1a631),
	.ram_block1a31(ram_block1a311),
	.address_reg_a_0(address_reg_a_0),
	.l1_w16_n0_mux_dataout(l1_w16_n0_mux_dataout1),
	.l1_w17_n0_mux_dataout(l1_w17_n0_mux_dataout1),
	.l1_w18_n0_mux_dataout(l1_w18_n0_mux_dataout1),
	.l1_w19_n0_mux_dataout(l1_w19_n0_mux_dataout1),
	.l1_w20_n0_mux_dataout(l1_w20_n0_mux_dataout1),
	.l1_w21_n0_mux_dataout(l1_w21_n0_mux_dataout1),
	.l1_w22_n0_mux_dataout(l1_w22_n0_mux_dataout1),
	.l1_w23_n0_mux_dataout(l1_w23_n0_mux_dataout1),
	.l1_w8_n0_mux_dataout(l1_w8_n0_mux_dataout1),
	.l1_w9_n0_mux_dataout(l1_w9_n0_mux_dataout1),
	.l1_w10_n0_mux_dataout(l1_w10_n0_mux_dataout1),
	.l1_w11_n0_mux_dataout(l1_w11_n0_mux_dataout1),
	.l1_w12_n0_mux_dataout(l1_w12_n0_mux_dataout1),
	.l1_w13_n0_mux_dataout(l1_w13_n0_mux_dataout1),
	.l1_w14_n0_mux_dataout(l1_w14_n0_mux_dataout1),
	.l1_w15_n0_mux_dataout(l1_w15_n0_mux_dataout1),
	.l1_w24_n0_mux_dataout(l1_w24_n0_mux_dataout1),
	.l1_w25_n0_mux_dataout(l1_w25_n0_mux_dataout1),
	.l1_w26_n0_mux_dataout(l1_w26_n0_mux_dataout1),
	.l1_w27_n0_mux_dataout(l1_w27_n0_mux_dataout1),
	.l1_w28_n0_mux_dataout(l1_w28_n0_mux_dataout1),
	.l1_w29_n0_mux_dataout(l1_w29_n0_mux_dataout1),
	.l1_w30_n0_mux_dataout(l1_w30_n0_mux_dataout1),
	.l1_w31_n0_mux_dataout(l1_w31_n0_mux_dataout1));

Computer_System_decode_5la_1 decode3(
	.eq_node_1(\decode3|eq_node[1]~0_combout ),
	.eq_node_0(\decode3|eq_node[0]~1_combout ),
	.onchip_sram_s2_address_13(address_b[13]),
	.onchip_sram_s2_chipselect(onchip_sram_s2_chipselect),
	.onchip_sram_s2_write(onchip_sram_s2_write));

Computer_System_decode_5la decode2(
	.readaddress_15(readaddress_15),
	.writeaddress_15(writeaddress_15),
	.saved_grant_0(saved_grant_0),
	.saved_grant_1(saved_grant_1),
	.wren(wren),
	.eq_node_1(\decode2|eq_node[1]~combout ),
	.eq_node_0(\decode2|eq_node[0]~combout ));

cyclonev_ram_block ram_block1a48(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a48_PORTADATAOUT_bus),
	.portbdataout(ram_block1a48_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena0";
defparam ram_block1a48.clk1_core_clock_enable = "ena1";
defparam ram_block1a48.clk1_input_clock_enable = "ena1";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a48.operation_mode = "bidir_dual_port";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 13;
defparam ram_block1a48.port_a_byte_enable_mask_width = 1;
defparam ram_block1a48.port_a_byte_size = 1;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "none";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 8192;
defparam ram_block1a48.port_a_first_bit_number = 16;
defparam ram_block1a48.port_a_last_address = 16383;
defparam ram_block1a48.port_a_logical_ram_depth = 16384;
defparam ram_block1a48.port_a_logical_ram_width = 32;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.port_b_address_clear = "none";
defparam ram_block1a48.port_b_address_clock = "clock1";
defparam ram_block1a48.port_b_address_width = 13;
defparam ram_block1a48.port_b_byte_enable_clock = "clock1";
defparam ram_block1a48.port_b_byte_enable_mask_width = 1;
defparam ram_block1a48.port_b_byte_size = 1;
defparam ram_block1a48.port_b_data_in_clock = "clock1";
defparam ram_block1a48.port_b_data_out_clear = "none";
defparam ram_block1a48.port_b_data_out_clock = "none";
defparam ram_block1a48.port_b_data_width = 1;
defparam ram_block1a48.port_b_first_address = 8192;
defparam ram_block1a48.port_b_first_bit_number = 16;
defparam ram_block1a48.port_b_last_address = 16383;
defparam ram_block1a48.port_b_logical_ram_depth = 16384;
defparam ram_block1a48.port_b_logical_ram_width = 32;
defparam ram_block1a48.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.port_b_read_enable_clock = "clock1";
defparam ram_block1a48.port_b_write_enable_clock = "clock1";
defparam ram_block1a48.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.clk1_input_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "bidir_dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 16384;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 13;
defparam ram_block1a16.port_b_byte_enable_clock = "clock1";
defparam ram_block1a16.port_b_byte_enable_mask_width = 1;
defparam ram_block1a16.port_b_byte_size = 1;
defparam ram_block1a16.port_b_data_in_clock = "clock1";
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 8191;
defparam ram_block1a16.port_b_logical_ram_depth = 16384;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.port_b_write_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a49(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a49_PORTADATAOUT_bus),
	.portbdataout(ram_block1a49_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena0";
defparam ram_block1a49.clk1_core_clock_enable = "ena1";
defparam ram_block1a49.clk1_input_clock_enable = "ena1";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a49.operation_mode = "bidir_dual_port";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 13;
defparam ram_block1a49.port_a_byte_enable_mask_width = 1;
defparam ram_block1a49.port_a_byte_size = 1;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "none";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 8192;
defparam ram_block1a49.port_a_first_bit_number = 17;
defparam ram_block1a49.port_a_last_address = 16383;
defparam ram_block1a49.port_a_logical_ram_depth = 16384;
defparam ram_block1a49.port_a_logical_ram_width = 32;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.port_b_address_clear = "none";
defparam ram_block1a49.port_b_address_clock = "clock1";
defparam ram_block1a49.port_b_address_width = 13;
defparam ram_block1a49.port_b_byte_enable_clock = "clock1";
defparam ram_block1a49.port_b_byte_enable_mask_width = 1;
defparam ram_block1a49.port_b_byte_size = 1;
defparam ram_block1a49.port_b_data_in_clock = "clock1";
defparam ram_block1a49.port_b_data_out_clear = "none";
defparam ram_block1a49.port_b_data_out_clock = "none";
defparam ram_block1a49.port_b_data_width = 1;
defparam ram_block1a49.port_b_first_address = 8192;
defparam ram_block1a49.port_b_first_bit_number = 17;
defparam ram_block1a49.port_b_last_address = 16383;
defparam ram_block1a49.port_b_logical_ram_depth = 16384;
defparam ram_block1a49.port_b_logical_ram_width = 32;
defparam ram_block1a49.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.port_b_read_enable_clock = "clock1";
defparam ram_block1a49.port_b_write_enable_clock = "clock1";
defparam ram_block1a49.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.clk1_input_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "bidir_dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 16384;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 13;
defparam ram_block1a17.port_b_byte_enable_clock = "clock1";
defparam ram_block1a17.port_b_byte_enable_mask_width = 1;
defparam ram_block1a17.port_b_byte_size = 1;
defparam ram_block1a17.port_b_data_in_clock = "clock1";
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 8191;
defparam ram_block1a17.port_b_logical_ram_depth = 16384;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.port_b_write_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a50(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a50_PORTADATAOUT_bus),
	.portbdataout(ram_block1a50_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena0";
defparam ram_block1a50.clk1_core_clock_enable = "ena1";
defparam ram_block1a50.clk1_input_clock_enable = "ena1";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a50.operation_mode = "bidir_dual_port";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 13;
defparam ram_block1a50.port_a_byte_enable_mask_width = 1;
defparam ram_block1a50.port_a_byte_size = 1;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "none";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 8192;
defparam ram_block1a50.port_a_first_bit_number = 18;
defparam ram_block1a50.port_a_last_address = 16383;
defparam ram_block1a50.port_a_logical_ram_depth = 16384;
defparam ram_block1a50.port_a_logical_ram_width = 32;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.port_b_address_clear = "none";
defparam ram_block1a50.port_b_address_clock = "clock1";
defparam ram_block1a50.port_b_address_width = 13;
defparam ram_block1a50.port_b_byte_enable_clock = "clock1";
defparam ram_block1a50.port_b_byte_enable_mask_width = 1;
defparam ram_block1a50.port_b_byte_size = 1;
defparam ram_block1a50.port_b_data_in_clock = "clock1";
defparam ram_block1a50.port_b_data_out_clear = "none";
defparam ram_block1a50.port_b_data_out_clock = "none";
defparam ram_block1a50.port_b_data_width = 1;
defparam ram_block1a50.port_b_first_address = 8192;
defparam ram_block1a50.port_b_first_bit_number = 18;
defparam ram_block1a50.port_b_last_address = 16383;
defparam ram_block1a50.port_b_logical_ram_depth = 16384;
defparam ram_block1a50.port_b_logical_ram_width = 32;
defparam ram_block1a50.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.port_b_read_enable_clock = "clock1";
defparam ram_block1a50.port_b_write_enable_clock = "clock1";
defparam ram_block1a50.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.clk1_input_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "bidir_dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 16384;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 13;
defparam ram_block1a18.port_b_byte_enable_clock = "clock1";
defparam ram_block1a18.port_b_byte_enable_mask_width = 1;
defparam ram_block1a18.port_b_byte_size = 1;
defparam ram_block1a18.port_b_data_in_clock = "clock1";
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 8191;
defparam ram_block1a18.port_b_logical_ram_depth = 16384;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.port_b_write_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a51(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a51_PORTADATAOUT_bus),
	.portbdataout(ram_block1a51_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena0";
defparam ram_block1a51.clk1_core_clock_enable = "ena1";
defparam ram_block1a51.clk1_input_clock_enable = "ena1";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a51.operation_mode = "bidir_dual_port";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 13;
defparam ram_block1a51.port_a_byte_enable_mask_width = 1;
defparam ram_block1a51.port_a_byte_size = 1;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "none";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 8192;
defparam ram_block1a51.port_a_first_bit_number = 19;
defparam ram_block1a51.port_a_last_address = 16383;
defparam ram_block1a51.port_a_logical_ram_depth = 16384;
defparam ram_block1a51.port_a_logical_ram_width = 32;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.port_b_address_clear = "none";
defparam ram_block1a51.port_b_address_clock = "clock1";
defparam ram_block1a51.port_b_address_width = 13;
defparam ram_block1a51.port_b_byte_enable_clock = "clock1";
defparam ram_block1a51.port_b_byte_enable_mask_width = 1;
defparam ram_block1a51.port_b_byte_size = 1;
defparam ram_block1a51.port_b_data_in_clock = "clock1";
defparam ram_block1a51.port_b_data_out_clear = "none";
defparam ram_block1a51.port_b_data_out_clock = "none";
defparam ram_block1a51.port_b_data_width = 1;
defparam ram_block1a51.port_b_first_address = 8192;
defparam ram_block1a51.port_b_first_bit_number = 19;
defparam ram_block1a51.port_b_last_address = 16383;
defparam ram_block1a51.port_b_logical_ram_depth = 16384;
defparam ram_block1a51.port_b_logical_ram_width = 32;
defparam ram_block1a51.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.port_b_read_enable_clock = "clock1";
defparam ram_block1a51.port_b_write_enable_clock = "clock1";
defparam ram_block1a51.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.clk1_input_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "bidir_dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 16384;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 13;
defparam ram_block1a19.port_b_byte_enable_clock = "clock1";
defparam ram_block1a19.port_b_byte_enable_mask_width = 1;
defparam ram_block1a19.port_b_byte_size = 1;
defparam ram_block1a19.port_b_data_in_clock = "clock1";
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 8191;
defparam ram_block1a19.port_b_logical_ram_depth = 16384;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.port_b_write_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a52(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a52_PORTADATAOUT_bus),
	.portbdataout(ram_block1a52_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena0";
defparam ram_block1a52.clk1_core_clock_enable = "ena1";
defparam ram_block1a52.clk1_input_clock_enable = "ena1";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a52.operation_mode = "bidir_dual_port";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 13;
defparam ram_block1a52.port_a_byte_enable_mask_width = 1;
defparam ram_block1a52.port_a_byte_size = 1;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "none";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 8192;
defparam ram_block1a52.port_a_first_bit_number = 20;
defparam ram_block1a52.port_a_last_address = 16383;
defparam ram_block1a52.port_a_logical_ram_depth = 16384;
defparam ram_block1a52.port_a_logical_ram_width = 32;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.port_b_address_clear = "none";
defparam ram_block1a52.port_b_address_clock = "clock1";
defparam ram_block1a52.port_b_address_width = 13;
defparam ram_block1a52.port_b_byte_enable_clock = "clock1";
defparam ram_block1a52.port_b_byte_enable_mask_width = 1;
defparam ram_block1a52.port_b_byte_size = 1;
defparam ram_block1a52.port_b_data_in_clock = "clock1";
defparam ram_block1a52.port_b_data_out_clear = "none";
defparam ram_block1a52.port_b_data_out_clock = "none";
defparam ram_block1a52.port_b_data_width = 1;
defparam ram_block1a52.port_b_first_address = 8192;
defparam ram_block1a52.port_b_first_bit_number = 20;
defparam ram_block1a52.port_b_last_address = 16383;
defparam ram_block1a52.port_b_logical_ram_depth = 16384;
defparam ram_block1a52.port_b_logical_ram_width = 32;
defparam ram_block1a52.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.port_b_read_enable_clock = "clock1";
defparam ram_block1a52.port_b_write_enable_clock = "clock1";
defparam ram_block1a52.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.clk1_input_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "bidir_dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 16384;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 13;
defparam ram_block1a20.port_b_byte_enable_clock = "clock1";
defparam ram_block1a20.port_b_byte_enable_mask_width = 1;
defparam ram_block1a20.port_b_byte_size = 1;
defparam ram_block1a20.port_b_data_in_clock = "clock1";
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 8191;
defparam ram_block1a20.port_b_logical_ram_depth = 16384;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.port_b_write_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a53(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a53_PORTADATAOUT_bus),
	.portbdataout(ram_block1a53_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena0";
defparam ram_block1a53.clk1_core_clock_enable = "ena1";
defparam ram_block1a53.clk1_input_clock_enable = "ena1";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a53.operation_mode = "bidir_dual_port";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 13;
defparam ram_block1a53.port_a_byte_enable_mask_width = 1;
defparam ram_block1a53.port_a_byte_size = 1;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "none";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 8192;
defparam ram_block1a53.port_a_first_bit_number = 21;
defparam ram_block1a53.port_a_last_address = 16383;
defparam ram_block1a53.port_a_logical_ram_depth = 16384;
defparam ram_block1a53.port_a_logical_ram_width = 32;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.port_b_address_clear = "none";
defparam ram_block1a53.port_b_address_clock = "clock1";
defparam ram_block1a53.port_b_address_width = 13;
defparam ram_block1a53.port_b_byte_enable_clock = "clock1";
defparam ram_block1a53.port_b_byte_enable_mask_width = 1;
defparam ram_block1a53.port_b_byte_size = 1;
defparam ram_block1a53.port_b_data_in_clock = "clock1";
defparam ram_block1a53.port_b_data_out_clear = "none";
defparam ram_block1a53.port_b_data_out_clock = "none";
defparam ram_block1a53.port_b_data_width = 1;
defparam ram_block1a53.port_b_first_address = 8192;
defparam ram_block1a53.port_b_first_bit_number = 21;
defparam ram_block1a53.port_b_last_address = 16383;
defparam ram_block1a53.port_b_logical_ram_depth = 16384;
defparam ram_block1a53.port_b_logical_ram_width = 32;
defparam ram_block1a53.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.port_b_read_enable_clock = "clock1";
defparam ram_block1a53.port_b_write_enable_clock = "clock1";
defparam ram_block1a53.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.clk1_input_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "bidir_dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 16384;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 13;
defparam ram_block1a21.port_b_byte_enable_clock = "clock1";
defparam ram_block1a21.port_b_byte_enable_mask_width = 1;
defparam ram_block1a21.port_b_byte_size = 1;
defparam ram_block1a21.port_b_data_in_clock = "clock1";
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 8191;
defparam ram_block1a21.port_b_logical_ram_depth = 16384;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.port_b_write_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a54(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a54_PORTADATAOUT_bus),
	.portbdataout(ram_block1a54_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena0";
defparam ram_block1a54.clk1_core_clock_enable = "ena1";
defparam ram_block1a54.clk1_input_clock_enable = "ena1";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a54.operation_mode = "bidir_dual_port";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 13;
defparam ram_block1a54.port_a_byte_enable_mask_width = 1;
defparam ram_block1a54.port_a_byte_size = 1;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "none";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 8192;
defparam ram_block1a54.port_a_first_bit_number = 22;
defparam ram_block1a54.port_a_last_address = 16383;
defparam ram_block1a54.port_a_logical_ram_depth = 16384;
defparam ram_block1a54.port_a_logical_ram_width = 32;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.port_b_address_clear = "none";
defparam ram_block1a54.port_b_address_clock = "clock1";
defparam ram_block1a54.port_b_address_width = 13;
defparam ram_block1a54.port_b_byte_enable_clock = "clock1";
defparam ram_block1a54.port_b_byte_enable_mask_width = 1;
defparam ram_block1a54.port_b_byte_size = 1;
defparam ram_block1a54.port_b_data_in_clock = "clock1";
defparam ram_block1a54.port_b_data_out_clear = "none";
defparam ram_block1a54.port_b_data_out_clock = "none";
defparam ram_block1a54.port_b_data_width = 1;
defparam ram_block1a54.port_b_first_address = 8192;
defparam ram_block1a54.port_b_first_bit_number = 22;
defparam ram_block1a54.port_b_last_address = 16383;
defparam ram_block1a54.port_b_logical_ram_depth = 16384;
defparam ram_block1a54.port_b_logical_ram_width = 32;
defparam ram_block1a54.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.port_b_read_enable_clock = "clock1";
defparam ram_block1a54.port_b_write_enable_clock = "clock1";
defparam ram_block1a54.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.clk1_input_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "bidir_dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 16384;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 13;
defparam ram_block1a22.port_b_byte_enable_clock = "clock1";
defparam ram_block1a22.port_b_byte_enable_mask_width = 1;
defparam ram_block1a22.port_b_byte_size = 1;
defparam ram_block1a22.port_b_data_in_clock = "clock1";
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 8191;
defparam ram_block1a22.port_b_logical_ram_depth = 16384;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.port_b_write_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a55(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a55_PORTADATAOUT_bus),
	.portbdataout(ram_block1a55_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena0";
defparam ram_block1a55.clk1_core_clock_enable = "ena1";
defparam ram_block1a55.clk1_input_clock_enable = "ena1";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a55.operation_mode = "bidir_dual_port";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 13;
defparam ram_block1a55.port_a_byte_enable_mask_width = 1;
defparam ram_block1a55.port_a_byte_size = 1;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "none";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 8192;
defparam ram_block1a55.port_a_first_bit_number = 23;
defparam ram_block1a55.port_a_last_address = 16383;
defparam ram_block1a55.port_a_logical_ram_depth = 16384;
defparam ram_block1a55.port_a_logical_ram_width = 32;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.port_b_address_clear = "none";
defparam ram_block1a55.port_b_address_clock = "clock1";
defparam ram_block1a55.port_b_address_width = 13;
defparam ram_block1a55.port_b_byte_enable_clock = "clock1";
defparam ram_block1a55.port_b_byte_enable_mask_width = 1;
defparam ram_block1a55.port_b_byte_size = 1;
defparam ram_block1a55.port_b_data_in_clock = "clock1";
defparam ram_block1a55.port_b_data_out_clear = "none";
defparam ram_block1a55.port_b_data_out_clock = "none";
defparam ram_block1a55.port_b_data_width = 1;
defparam ram_block1a55.port_b_first_address = 8192;
defparam ram_block1a55.port_b_first_bit_number = 23;
defparam ram_block1a55.port_b_last_address = 16383;
defparam ram_block1a55.port_b_logical_ram_depth = 16384;
defparam ram_block1a55.port_b_logical_ram_width = 32;
defparam ram_block1a55.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.port_b_read_enable_clock = "clock1";
defparam ram_block1a55.port_b_write_enable_clock = "clock1";
defparam ram_block1a55.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.clk1_input_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "bidir_dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 16384;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 13;
defparam ram_block1a23.port_b_byte_enable_clock = "clock1";
defparam ram_block1a23.port_b_byte_enable_mask_width = 1;
defparam ram_block1a23.port_b_byte_size = 1;
defparam ram_block1a23.port_b_data_in_clock = "clock1";
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 8191;
defparam ram_block1a23.port_b_logical_ram_depth = 16384;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.port_b_write_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(address_b[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken1),
	.q(\address_reg_b[0]~q ),
	.prn(vcc));
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";

cyclonev_ram_block ram_block1a32(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a32_PORTADATAOUT_bus),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena0";
defparam ram_block1a32.clk1_core_clock_enable = "ena1";
defparam ram_block1a32.clk1_input_clock_enable = "ena1";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "bidir_dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 13;
defparam ram_block1a32.port_a_byte_enable_mask_width = 1;
defparam ram_block1a32.port_a_byte_size = 1;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 8192;
defparam ram_block1a32.port_a_first_bit_number = 0;
defparam ram_block1a32.port_a_last_address = 16383;
defparam ram_block1a32.port_a_logical_ram_depth = 16384;
defparam ram_block1a32.port_a_logical_ram_width = 32;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 13;
defparam ram_block1a32.port_b_byte_enable_clock = "clock1";
defparam ram_block1a32.port_b_byte_enable_mask_width = 1;
defparam ram_block1a32.port_b_byte_size = 1;
defparam ram_block1a32.port_b_data_in_clock = "clock1";
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "none";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 8192;
defparam ram_block1a32.port_b_first_bit_number = 0;
defparam ram_block1a32.port_b_last_address = 16383;
defparam ram_block1a32.port_b_logical_ram_depth = 16384;
defparam ram_block1a32.port_b_logical_ram_width = 32;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.port_b_write_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 16384;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 13;
defparam ram_block1a0.port_b_byte_enable_clock = "clock1";
defparam ram_block1a0.port_b_byte_enable_mask_width = 1;
defparam ram_block1a0.port_b_byte_size = 1;
defparam ram_block1a0.port_b_data_in_clock = "clock1";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 8191;
defparam ram_block1a0.port_b_logical_ram_depth = 16384;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.port_b_write_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a33(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a33_PORTADATAOUT_bus),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena0";
defparam ram_block1a33.clk1_core_clock_enable = "ena1";
defparam ram_block1a33.clk1_input_clock_enable = "ena1";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "bidir_dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 13;
defparam ram_block1a33.port_a_byte_enable_mask_width = 1;
defparam ram_block1a33.port_a_byte_size = 1;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 8192;
defparam ram_block1a33.port_a_first_bit_number = 1;
defparam ram_block1a33.port_a_last_address = 16383;
defparam ram_block1a33.port_a_logical_ram_depth = 16384;
defparam ram_block1a33.port_a_logical_ram_width = 32;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 13;
defparam ram_block1a33.port_b_byte_enable_clock = "clock1";
defparam ram_block1a33.port_b_byte_enable_mask_width = 1;
defparam ram_block1a33.port_b_byte_size = 1;
defparam ram_block1a33.port_b_data_in_clock = "clock1";
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "none";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 8192;
defparam ram_block1a33.port_b_first_bit_number = 1;
defparam ram_block1a33.port_b_last_address = 16383;
defparam ram_block1a33.port_b_logical_ram_depth = 16384;
defparam ram_block1a33.port_b_logical_ram_width = 32;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.port_b_write_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 16384;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 13;
defparam ram_block1a1.port_b_byte_enable_clock = "clock1";
defparam ram_block1a1.port_b_byte_enable_mask_width = 1;
defparam ram_block1a1.port_b_byte_size = 1;
defparam ram_block1a1.port_b_data_in_clock = "clock1";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 8191;
defparam ram_block1a1.port_b_logical_ram_depth = 16384;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.port_b_write_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a34(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a34_PORTADATAOUT_bus),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena0";
defparam ram_block1a34.clk1_core_clock_enable = "ena1";
defparam ram_block1a34.clk1_input_clock_enable = "ena1";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "bidir_dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 13;
defparam ram_block1a34.port_a_byte_enable_mask_width = 1;
defparam ram_block1a34.port_a_byte_size = 1;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 8192;
defparam ram_block1a34.port_a_first_bit_number = 2;
defparam ram_block1a34.port_a_last_address = 16383;
defparam ram_block1a34.port_a_logical_ram_depth = 16384;
defparam ram_block1a34.port_a_logical_ram_width = 32;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 13;
defparam ram_block1a34.port_b_byte_enable_clock = "clock1";
defparam ram_block1a34.port_b_byte_enable_mask_width = 1;
defparam ram_block1a34.port_b_byte_size = 1;
defparam ram_block1a34.port_b_data_in_clock = "clock1";
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "none";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 8192;
defparam ram_block1a34.port_b_first_bit_number = 2;
defparam ram_block1a34.port_b_last_address = 16383;
defparam ram_block1a34.port_b_logical_ram_depth = 16384;
defparam ram_block1a34.port_b_logical_ram_width = 32;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.port_b_write_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 16384;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 13;
defparam ram_block1a2.port_b_byte_enable_clock = "clock1";
defparam ram_block1a2.port_b_byte_enable_mask_width = 1;
defparam ram_block1a2.port_b_byte_size = 1;
defparam ram_block1a2.port_b_data_in_clock = "clock1";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 8191;
defparam ram_block1a2.port_b_logical_ram_depth = 16384;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.port_b_write_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a35(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a35_PORTADATAOUT_bus),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena0";
defparam ram_block1a35.clk1_core_clock_enable = "ena1";
defparam ram_block1a35.clk1_input_clock_enable = "ena1";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "bidir_dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 13;
defparam ram_block1a35.port_a_byte_enable_mask_width = 1;
defparam ram_block1a35.port_a_byte_size = 1;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 8192;
defparam ram_block1a35.port_a_first_bit_number = 3;
defparam ram_block1a35.port_a_last_address = 16383;
defparam ram_block1a35.port_a_logical_ram_depth = 16384;
defparam ram_block1a35.port_a_logical_ram_width = 32;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 13;
defparam ram_block1a35.port_b_byte_enable_clock = "clock1";
defparam ram_block1a35.port_b_byte_enable_mask_width = 1;
defparam ram_block1a35.port_b_byte_size = 1;
defparam ram_block1a35.port_b_data_in_clock = "clock1";
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "none";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 8192;
defparam ram_block1a35.port_b_first_bit_number = 3;
defparam ram_block1a35.port_b_last_address = 16383;
defparam ram_block1a35.port_b_logical_ram_depth = 16384;
defparam ram_block1a35.port_b_logical_ram_width = 32;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.port_b_write_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 16384;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 13;
defparam ram_block1a3.port_b_byte_enable_clock = "clock1";
defparam ram_block1a3.port_b_byte_enable_mask_width = 1;
defparam ram_block1a3.port_b_byte_size = 1;
defparam ram_block1a3.port_b_data_in_clock = "clock1";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 8191;
defparam ram_block1a3.port_b_logical_ram_depth = 16384;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.port_b_write_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a36(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a36_PORTADATAOUT_bus),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena0";
defparam ram_block1a36.clk1_core_clock_enable = "ena1";
defparam ram_block1a36.clk1_input_clock_enable = "ena1";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "bidir_dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 13;
defparam ram_block1a36.port_a_byte_enable_mask_width = 1;
defparam ram_block1a36.port_a_byte_size = 1;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 8192;
defparam ram_block1a36.port_a_first_bit_number = 4;
defparam ram_block1a36.port_a_last_address = 16383;
defparam ram_block1a36.port_a_logical_ram_depth = 16384;
defparam ram_block1a36.port_a_logical_ram_width = 32;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 13;
defparam ram_block1a36.port_b_byte_enable_clock = "clock1";
defparam ram_block1a36.port_b_byte_enable_mask_width = 1;
defparam ram_block1a36.port_b_byte_size = 1;
defparam ram_block1a36.port_b_data_in_clock = "clock1";
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "none";
defparam ram_block1a36.port_b_data_width = 1;
defparam ram_block1a36.port_b_first_address = 8192;
defparam ram_block1a36.port_b_first_bit_number = 4;
defparam ram_block1a36.port_b_last_address = 16383;
defparam ram_block1a36.port_b_logical_ram_depth = 16384;
defparam ram_block1a36.port_b_logical_ram_width = 32;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.port_b_write_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 16384;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 13;
defparam ram_block1a4.port_b_byte_enable_clock = "clock1";
defparam ram_block1a4.port_b_byte_enable_mask_width = 1;
defparam ram_block1a4.port_b_byte_size = 1;
defparam ram_block1a4.port_b_data_in_clock = "clock1";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 8191;
defparam ram_block1a4.port_b_logical_ram_depth = 16384;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.port_b_write_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a37(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a37_PORTADATAOUT_bus),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena0";
defparam ram_block1a37.clk1_core_clock_enable = "ena1";
defparam ram_block1a37.clk1_input_clock_enable = "ena1";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "bidir_dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 13;
defparam ram_block1a37.port_a_byte_enable_mask_width = 1;
defparam ram_block1a37.port_a_byte_size = 1;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 8192;
defparam ram_block1a37.port_a_first_bit_number = 5;
defparam ram_block1a37.port_a_last_address = 16383;
defparam ram_block1a37.port_a_logical_ram_depth = 16384;
defparam ram_block1a37.port_a_logical_ram_width = 32;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 13;
defparam ram_block1a37.port_b_byte_enable_clock = "clock1";
defparam ram_block1a37.port_b_byte_enable_mask_width = 1;
defparam ram_block1a37.port_b_byte_size = 1;
defparam ram_block1a37.port_b_data_in_clock = "clock1";
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "none";
defparam ram_block1a37.port_b_data_width = 1;
defparam ram_block1a37.port_b_first_address = 8192;
defparam ram_block1a37.port_b_first_bit_number = 5;
defparam ram_block1a37.port_b_last_address = 16383;
defparam ram_block1a37.port_b_logical_ram_depth = 16384;
defparam ram_block1a37.port_b_logical_ram_width = 32;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.port_b_write_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 16384;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 13;
defparam ram_block1a5.port_b_byte_enable_clock = "clock1";
defparam ram_block1a5.port_b_byte_enable_mask_width = 1;
defparam ram_block1a5.port_b_byte_size = 1;
defparam ram_block1a5.port_b_data_in_clock = "clock1";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 8191;
defparam ram_block1a5.port_b_logical_ram_depth = 16384;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.port_b_write_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a38(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a38_PORTADATAOUT_bus),
	.portbdataout(ram_block1a38_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena0";
defparam ram_block1a38.clk1_core_clock_enable = "ena1";
defparam ram_block1a38.clk1_input_clock_enable = "ena1";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a38.operation_mode = "bidir_dual_port";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 13;
defparam ram_block1a38.port_a_byte_enable_mask_width = 1;
defparam ram_block1a38.port_a_byte_size = 1;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "none";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 8192;
defparam ram_block1a38.port_a_first_bit_number = 6;
defparam ram_block1a38.port_a_last_address = 16383;
defparam ram_block1a38.port_a_logical_ram_depth = 16384;
defparam ram_block1a38.port_a_logical_ram_width = 32;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.port_b_address_clear = "none";
defparam ram_block1a38.port_b_address_clock = "clock1";
defparam ram_block1a38.port_b_address_width = 13;
defparam ram_block1a38.port_b_byte_enable_clock = "clock1";
defparam ram_block1a38.port_b_byte_enable_mask_width = 1;
defparam ram_block1a38.port_b_byte_size = 1;
defparam ram_block1a38.port_b_data_in_clock = "clock1";
defparam ram_block1a38.port_b_data_out_clear = "none";
defparam ram_block1a38.port_b_data_out_clock = "none";
defparam ram_block1a38.port_b_data_width = 1;
defparam ram_block1a38.port_b_first_address = 8192;
defparam ram_block1a38.port_b_first_bit_number = 6;
defparam ram_block1a38.port_b_last_address = 16383;
defparam ram_block1a38.port_b_logical_ram_depth = 16384;
defparam ram_block1a38.port_b_logical_ram_width = 32;
defparam ram_block1a38.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.port_b_read_enable_clock = "clock1";
defparam ram_block1a38.port_b_write_enable_clock = "clock1";
defparam ram_block1a38.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 16384;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 13;
defparam ram_block1a6.port_b_byte_enable_clock = "clock1";
defparam ram_block1a6.port_b_byte_enable_mask_width = 1;
defparam ram_block1a6.port_b_byte_size = 1;
defparam ram_block1a6.port_b_data_in_clock = "clock1";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 8191;
defparam ram_block1a6.port_b_logical_ram_depth = 16384;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.port_b_write_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a39(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a39_PORTADATAOUT_bus),
	.portbdataout(ram_block1a39_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena0";
defparam ram_block1a39.clk1_core_clock_enable = "ena1";
defparam ram_block1a39.clk1_input_clock_enable = "ena1";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a39.operation_mode = "bidir_dual_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 13;
defparam ram_block1a39.port_a_byte_enable_mask_width = 1;
defparam ram_block1a39.port_a_byte_size = 1;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 8192;
defparam ram_block1a39.port_a_first_bit_number = 7;
defparam ram_block1a39.port_a_last_address = 16383;
defparam ram_block1a39.port_a_logical_ram_depth = 16384;
defparam ram_block1a39.port_a_logical_ram_width = 32;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_address_clear = "none";
defparam ram_block1a39.port_b_address_clock = "clock1";
defparam ram_block1a39.port_b_address_width = 13;
defparam ram_block1a39.port_b_byte_enable_clock = "clock1";
defparam ram_block1a39.port_b_byte_enable_mask_width = 1;
defparam ram_block1a39.port_b_byte_size = 1;
defparam ram_block1a39.port_b_data_in_clock = "clock1";
defparam ram_block1a39.port_b_data_out_clear = "none";
defparam ram_block1a39.port_b_data_out_clock = "none";
defparam ram_block1a39.port_b_data_width = 1;
defparam ram_block1a39.port_b_first_address = 8192;
defparam ram_block1a39.port_b_first_bit_number = 7;
defparam ram_block1a39.port_b_last_address = 16383;
defparam ram_block1a39.port_b_logical_ram_depth = 16384;
defparam ram_block1a39.port_b_logical_ram_width = 32;
defparam ram_block1a39.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_read_enable_clock = "clock1";
defparam ram_block1a39.port_b_write_enable_clock = "clock1";
defparam ram_block1a39.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 16384;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 13;
defparam ram_block1a7.port_b_byte_enable_clock = "clock1";
defparam ram_block1a7.port_b_byte_enable_mask_width = 1;
defparam ram_block1a7.port_b_byte_size = 1;
defparam ram_block1a7.port_b_data_in_clock = "clock1";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 8191;
defparam ram_block1a7.port_b_logical_ram_depth = 16384;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.port_b_write_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a40(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a40_PORTADATAOUT_bus),
	.portbdataout(ram_block1a40_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena0";
defparam ram_block1a40.clk1_core_clock_enable = "ena1";
defparam ram_block1a40.clk1_input_clock_enable = "ena1";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a40.operation_mode = "bidir_dual_port";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 13;
defparam ram_block1a40.port_a_byte_enable_mask_width = 1;
defparam ram_block1a40.port_a_byte_size = 1;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "none";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 8192;
defparam ram_block1a40.port_a_first_bit_number = 8;
defparam ram_block1a40.port_a_last_address = 16383;
defparam ram_block1a40.port_a_logical_ram_depth = 16384;
defparam ram_block1a40.port_a_logical_ram_width = 32;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.port_b_address_clear = "none";
defparam ram_block1a40.port_b_address_clock = "clock1";
defparam ram_block1a40.port_b_address_width = 13;
defparam ram_block1a40.port_b_byte_enable_clock = "clock1";
defparam ram_block1a40.port_b_byte_enable_mask_width = 1;
defparam ram_block1a40.port_b_byte_size = 1;
defparam ram_block1a40.port_b_data_in_clock = "clock1";
defparam ram_block1a40.port_b_data_out_clear = "none";
defparam ram_block1a40.port_b_data_out_clock = "none";
defparam ram_block1a40.port_b_data_width = 1;
defparam ram_block1a40.port_b_first_address = 8192;
defparam ram_block1a40.port_b_first_bit_number = 8;
defparam ram_block1a40.port_b_last_address = 16383;
defparam ram_block1a40.port_b_logical_ram_depth = 16384;
defparam ram_block1a40.port_b_logical_ram_width = 32;
defparam ram_block1a40.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.port_b_read_enable_clock = "clock1";
defparam ram_block1a40.port_b_write_enable_clock = "clock1";
defparam ram_block1a40.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 16384;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 13;
defparam ram_block1a8.port_b_byte_enable_clock = "clock1";
defparam ram_block1a8.port_b_byte_enable_mask_width = 1;
defparam ram_block1a8.port_b_byte_size = 1;
defparam ram_block1a8.port_b_data_in_clock = "clock1";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 8191;
defparam ram_block1a8.port_b_logical_ram_depth = 16384;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.port_b_write_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a41(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a41_PORTADATAOUT_bus),
	.portbdataout(ram_block1a41_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena0";
defparam ram_block1a41.clk1_core_clock_enable = "ena1";
defparam ram_block1a41.clk1_input_clock_enable = "ena1";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a41.operation_mode = "bidir_dual_port";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 13;
defparam ram_block1a41.port_a_byte_enable_mask_width = 1;
defparam ram_block1a41.port_a_byte_size = 1;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "none";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 8192;
defparam ram_block1a41.port_a_first_bit_number = 9;
defparam ram_block1a41.port_a_last_address = 16383;
defparam ram_block1a41.port_a_logical_ram_depth = 16384;
defparam ram_block1a41.port_a_logical_ram_width = 32;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.port_b_address_clear = "none";
defparam ram_block1a41.port_b_address_clock = "clock1";
defparam ram_block1a41.port_b_address_width = 13;
defparam ram_block1a41.port_b_byte_enable_clock = "clock1";
defparam ram_block1a41.port_b_byte_enable_mask_width = 1;
defparam ram_block1a41.port_b_byte_size = 1;
defparam ram_block1a41.port_b_data_in_clock = "clock1";
defparam ram_block1a41.port_b_data_out_clear = "none";
defparam ram_block1a41.port_b_data_out_clock = "none";
defparam ram_block1a41.port_b_data_width = 1;
defparam ram_block1a41.port_b_first_address = 8192;
defparam ram_block1a41.port_b_first_bit_number = 9;
defparam ram_block1a41.port_b_last_address = 16383;
defparam ram_block1a41.port_b_logical_ram_depth = 16384;
defparam ram_block1a41.port_b_logical_ram_width = 32;
defparam ram_block1a41.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.port_b_read_enable_clock = "clock1";
defparam ram_block1a41.port_b_write_enable_clock = "clock1";
defparam ram_block1a41.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 16384;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 13;
defparam ram_block1a9.port_b_byte_enable_clock = "clock1";
defparam ram_block1a9.port_b_byte_enable_mask_width = 1;
defparam ram_block1a9.port_b_byte_size = 1;
defparam ram_block1a9.port_b_data_in_clock = "clock1";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 8191;
defparam ram_block1a9.port_b_logical_ram_depth = 16384;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.port_b_write_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a42(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a42_PORTADATAOUT_bus),
	.portbdataout(ram_block1a42_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena0";
defparam ram_block1a42.clk1_core_clock_enable = "ena1";
defparam ram_block1a42.clk1_input_clock_enable = "ena1";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a42.operation_mode = "bidir_dual_port";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 13;
defparam ram_block1a42.port_a_byte_enable_mask_width = 1;
defparam ram_block1a42.port_a_byte_size = 1;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "none";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 8192;
defparam ram_block1a42.port_a_first_bit_number = 10;
defparam ram_block1a42.port_a_last_address = 16383;
defparam ram_block1a42.port_a_logical_ram_depth = 16384;
defparam ram_block1a42.port_a_logical_ram_width = 32;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.port_b_address_clear = "none";
defparam ram_block1a42.port_b_address_clock = "clock1";
defparam ram_block1a42.port_b_address_width = 13;
defparam ram_block1a42.port_b_byte_enable_clock = "clock1";
defparam ram_block1a42.port_b_byte_enable_mask_width = 1;
defparam ram_block1a42.port_b_byte_size = 1;
defparam ram_block1a42.port_b_data_in_clock = "clock1";
defparam ram_block1a42.port_b_data_out_clear = "none";
defparam ram_block1a42.port_b_data_out_clock = "none";
defparam ram_block1a42.port_b_data_width = 1;
defparam ram_block1a42.port_b_first_address = 8192;
defparam ram_block1a42.port_b_first_bit_number = 10;
defparam ram_block1a42.port_b_last_address = 16383;
defparam ram_block1a42.port_b_logical_ram_depth = 16384;
defparam ram_block1a42.port_b_logical_ram_width = 32;
defparam ram_block1a42.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.port_b_read_enable_clock = "clock1";
defparam ram_block1a42.port_b_write_enable_clock = "clock1";
defparam ram_block1a42.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 16384;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 13;
defparam ram_block1a10.port_b_byte_enable_clock = "clock1";
defparam ram_block1a10.port_b_byte_enable_mask_width = 1;
defparam ram_block1a10.port_b_byte_size = 1;
defparam ram_block1a10.port_b_data_in_clock = "clock1";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 8191;
defparam ram_block1a10.port_b_logical_ram_depth = 16384;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.port_b_write_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a43(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a43_PORTADATAOUT_bus),
	.portbdataout(ram_block1a43_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena0";
defparam ram_block1a43.clk1_core_clock_enable = "ena1";
defparam ram_block1a43.clk1_input_clock_enable = "ena1";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a43.operation_mode = "bidir_dual_port";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 13;
defparam ram_block1a43.port_a_byte_enable_mask_width = 1;
defparam ram_block1a43.port_a_byte_size = 1;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "none";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 8192;
defparam ram_block1a43.port_a_first_bit_number = 11;
defparam ram_block1a43.port_a_last_address = 16383;
defparam ram_block1a43.port_a_logical_ram_depth = 16384;
defparam ram_block1a43.port_a_logical_ram_width = 32;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.port_b_address_clear = "none";
defparam ram_block1a43.port_b_address_clock = "clock1";
defparam ram_block1a43.port_b_address_width = 13;
defparam ram_block1a43.port_b_byte_enable_clock = "clock1";
defparam ram_block1a43.port_b_byte_enable_mask_width = 1;
defparam ram_block1a43.port_b_byte_size = 1;
defparam ram_block1a43.port_b_data_in_clock = "clock1";
defparam ram_block1a43.port_b_data_out_clear = "none";
defparam ram_block1a43.port_b_data_out_clock = "none";
defparam ram_block1a43.port_b_data_width = 1;
defparam ram_block1a43.port_b_first_address = 8192;
defparam ram_block1a43.port_b_first_bit_number = 11;
defparam ram_block1a43.port_b_last_address = 16383;
defparam ram_block1a43.port_b_logical_ram_depth = 16384;
defparam ram_block1a43.port_b_logical_ram_width = 32;
defparam ram_block1a43.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.port_b_read_enable_clock = "clock1";
defparam ram_block1a43.port_b_write_enable_clock = "clock1";
defparam ram_block1a43.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 16384;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 13;
defparam ram_block1a11.port_b_byte_enable_clock = "clock1";
defparam ram_block1a11.port_b_byte_enable_mask_width = 1;
defparam ram_block1a11.port_b_byte_size = 1;
defparam ram_block1a11.port_b_data_in_clock = "clock1";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 8191;
defparam ram_block1a11.port_b_logical_ram_depth = 16384;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.port_b_write_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a44(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a44_PORTADATAOUT_bus),
	.portbdataout(ram_block1a44_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena0";
defparam ram_block1a44.clk1_core_clock_enable = "ena1";
defparam ram_block1a44.clk1_input_clock_enable = "ena1";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a44.operation_mode = "bidir_dual_port";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 13;
defparam ram_block1a44.port_a_byte_enable_mask_width = 1;
defparam ram_block1a44.port_a_byte_size = 1;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "none";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 8192;
defparam ram_block1a44.port_a_first_bit_number = 12;
defparam ram_block1a44.port_a_last_address = 16383;
defparam ram_block1a44.port_a_logical_ram_depth = 16384;
defparam ram_block1a44.port_a_logical_ram_width = 32;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.port_b_address_clear = "none";
defparam ram_block1a44.port_b_address_clock = "clock1";
defparam ram_block1a44.port_b_address_width = 13;
defparam ram_block1a44.port_b_byte_enable_clock = "clock1";
defparam ram_block1a44.port_b_byte_enable_mask_width = 1;
defparam ram_block1a44.port_b_byte_size = 1;
defparam ram_block1a44.port_b_data_in_clock = "clock1";
defparam ram_block1a44.port_b_data_out_clear = "none";
defparam ram_block1a44.port_b_data_out_clock = "none";
defparam ram_block1a44.port_b_data_width = 1;
defparam ram_block1a44.port_b_first_address = 8192;
defparam ram_block1a44.port_b_first_bit_number = 12;
defparam ram_block1a44.port_b_last_address = 16383;
defparam ram_block1a44.port_b_logical_ram_depth = 16384;
defparam ram_block1a44.port_b_logical_ram_width = 32;
defparam ram_block1a44.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.port_b_read_enable_clock = "clock1";
defparam ram_block1a44.port_b_write_enable_clock = "clock1";
defparam ram_block1a44.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 16384;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 13;
defparam ram_block1a12.port_b_byte_enable_clock = "clock1";
defparam ram_block1a12.port_b_byte_enable_mask_width = 1;
defparam ram_block1a12.port_b_byte_size = 1;
defparam ram_block1a12.port_b_data_in_clock = "clock1";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 8191;
defparam ram_block1a12.port_b_logical_ram_depth = 16384;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.port_b_write_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a45(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a45_PORTADATAOUT_bus),
	.portbdataout(ram_block1a45_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena0";
defparam ram_block1a45.clk1_core_clock_enable = "ena1";
defparam ram_block1a45.clk1_input_clock_enable = "ena1";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a45.operation_mode = "bidir_dual_port";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 13;
defparam ram_block1a45.port_a_byte_enable_mask_width = 1;
defparam ram_block1a45.port_a_byte_size = 1;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "none";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 8192;
defparam ram_block1a45.port_a_first_bit_number = 13;
defparam ram_block1a45.port_a_last_address = 16383;
defparam ram_block1a45.port_a_logical_ram_depth = 16384;
defparam ram_block1a45.port_a_logical_ram_width = 32;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.port_b_address_clear = "none";
defparam ram_block1a45.port_b_address_clock = "clock1";
defparam ram_block1a45.port_b_address_width = 13;
defparam ram_block1a45.port_b_byte_enable_clock = "clock1";
defparam ram_block1a45.port_b_byte_enable_mask_width = 1;
defparam ram_block1a45.port_b_byte_size = 1;
defparam ram_block1a45.port_b_data_in_clock = "clock1";
defparam ram_block1a45.port_b_data_out_clear = "none";
defparam ram_block1a45.port_b_data_out_clock = "none";
defparam ram_block1a45.port_b_data_width = 1;
defparam ram_block1a45.port_b_first_address = 8192;
defparam ram_block1a45.port_b_first_bit_number = 13;
defparam ram_block1a45.port_b_last_address = 16383;
defparam ram_block1a45.port_b_logical_ram_depth = 16384;
defparam ram_block1a45.port_b_logical_ram_width = 32;
defparam ram_block1a45.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.port_b_read_enable_clock = "clock1";
defparam ram_block1a45.port_b_write_enable_clock = "clock1";
defparam ram_block1a45.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 16384;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 13;
defparam ram_block1a13.port_b_byte_enable_clock = "clock1";
defparam ram_block1a13.port_b_byte_enable_mask_width = 1;
defparam ram_block1a13.port_b_byte_size = 1;
defparam ram_block1a13.port_b_data_in_clock = "clock1";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 8191;
defparam ram_block1a13.port_b_logical_ram_depth = 16384;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.port_b_write_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a46(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a46_PORTADATAOUT_bus),
	.portbdataout(ram_block1a46_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena0";
defparam ram_block1a46.clk1_core_clock_enable = "ena1";
defparam ram_block1a46.clk1_input_clock_enable = "ena1";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a46.operation_mode = "bidir_dual_port";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 13;
defparam ram_block1a46.port_a_byte_enable_mask_width = 1;
defparam ram_block1a46.port_a_byte_size = 1;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "none";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 8192;
defparam ram_block1a46.port_a_first_bit_number = 14;
defparam ram_block1a46.port_a_last_address = 16383;
defparam ram_block1a46.port_a_logical_ram_depth = 16384;
defparam ram_block1a46.port_a_logical_ram_width = 32;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.port_b_address_clear = "none";
defparam ram_block1a46.port_b_address_clock = "clock1";
defparam ram_block1a46.port_b_address_width = 13;
defparam ram_block1a46.port_b_byte_enable_clock = "clock1";
defparam ram_block1a46.port_b_byte_enable_mask_width = 1;
defparam ram_block1a46.port_b_byte_size = 1;
defparam ram_block1a46.port_b_data_in_clock = "clock1";
defparam ram_block1a46.port_b_data_out_clear = "none";
defparam ram_block1a46.port_b_data_out_clock = "none";
defparam ram_block1a46.port_b_data_width = 1;
defparam ram_block1a46.port_b_first_address = 8192;
defparam ram_block1a46.port_b_first_bit_number = 14;
defparam ram_block1a46.port_b_last_address = 16383;
defparam ram_block1a46.port_b_logical_ram_depth = 16384;
defparam ram_block1a46.port_b_logical_ram_width = 32;
defparam ram_block1a46.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.port_b_read_enable_clock = "clock1";
defparam ram_block1a46.port_b_write_enable_clock = "clock1";
defparam ram_block1a46.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 16384;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 13;
defparam ram_block1a14.port_b_byte_enable_clock = "clock1";
defparam ram_block1a14.port_b_byte_enable_mask_width = 1;
defparam ram_block1a14.port_b_byte_size = 1;
defparam ram_block1a14.port_b_data_in_clock = "clock1";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 8191;
defparam ram_block1a14.port_b_logical_ram_depth = 16384;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.port_b_write_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a47(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a47_PORTADATAOUT_bus),
	.portbdataout(ram_block1a47_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena0";
defparam ram_block1a47.clk1_core_clock_enable = "ena1";
defparam ram_block1a47.clk1_input_clock_enable = "ena1";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a47.operation_mode = "bidir_dual_port";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 13;
defparam ram_block1a47.port_a_byte_enable_mask_width = 1;
defparam ram_block1a47.port_a_byte_size = 1;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "none";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 8192;
defparam ram_block1a47.port_a_first_bit_number = 15;
defparam ram_block1a47.port_a_last_address = 16383;
defparam ram_block1a47.port_a_logical_ram_depth = 16384;
defparam ram_block1a47.port_a_logical_ram_width = 32;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.port_b_address_clear = "none";
defparam ram_block1a47.port_b_address_clock = "clock1";
defparam ram_block1a47.port_b_address_width = 13;
defparam ram_block1a47.port_b_byte_enable_clock = "clock1";
defparam ram_block1a47.port_b_byte_enable_mask_width = 1;
defparam ram_block1a47.port_b_byte_size = 1;
defparam ram_block1a47.port_b_data_in_clock = "clock1";
defparam ram_block1a47.port_b_data_out_clear = "none";
defparam ram_block1a47.port_b_data_out_clock = "none";
defparam ram_block1a47.port_b_data_width = 1;
defparam ram_block1a47.port_b_first_address = 8192;
defparam ram_block1a47.port_b_first_bit_number = 15;
defparam ram_block1a47.port_b_last_address = 16383;
defparam ram_block1a47.port_b_logical_ram_depth = 16384;
defparam ram_block1a47.port_b_logical_ram_width = 32;
defparam ram_block1a47.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.port_b_read_enable_clock = "clock1";
defparam ram_block1a47.port_b_write_enable_clock = "clock1";
defparam ram_block1a47.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 16384;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 13;
defparam ram_block1a15.port_b_byte_enable_clock = "clock1";
defparam ram_block1a15.port_b_byte_enable_mask_width = 1;
defparam ram_block1a15.port_b_byte_size = 1;
defparam ram_block1a15.port_b_data_in_clock = "clock1";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 8191;
defparam ram_block1a15.port_b_logical_ram_depth = 16384;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.port_b_write_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a56(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a56_PORTADATAOUT_bus),
	.portbdataout(ram_block1a56_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena0";
defparam ram_block1a56.clk1_core_clock_enable = "ena1";
defparam ram_block1a56.clk1_input_clock_enable = "ena1";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a56.operation_mode = "bidir_dual_port";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 13;
defparam ram_block1a56.port_a_byte_enable_mask_width = 1;
defparam ram_block1a56.port_a_byte_size = 1;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "none";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 8192;
defparam ram_block1a56.port_a_first_bit_number = 24;
defparam ram_block1a56.port_a_last_address = 16383;
defparam ram_block1a56.port_a_logical_ram_depth = 16384;
defparam ram_block1a56.port_a_logical_ram_width = 32;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.port_b_address_clear = "none";
defparam ram_block1a56.port_b_address_clock = "clock1";
defparam ram_block1a56.port_b_address_width = 13;
defparam ram_block1a56.port_b_byte_enable_clock = "clock1";
defparam ram_block1a56.port_b_byte_enable_mask_width = 1;
defparam ram_block1a56.port_b_byte_size = 1;
defparam ram_block1a56.port_b_data_in_clock = "clock1";
defparam ram_block1a56.port_b_data_out_clear = "none";
defparam ram_block1a56.port_b_data_out_clock = "none";
defparam ram_block1a56.port_b_data_width = 1;
defparam ram_block1a56.port_b_first_address = 8192;
defparam ram_block1a56.port_b_first_bit_number = 24;
defparam ram_block1a56.port_b_last_address = 16383;
defparam ram_block1a56.port_b_logical_ram_depth = 16384;
defparam ram_block1a56.port_b_logical_ram_width = 32;
defparam ram_block1a56.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.port_b_read_enable_clock = "clock1";
defparam ram_block1a56.port_b_write_enable_clock = "clock1";
defparam ram_block1a56.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.clk1_input_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "bidir_dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 16384;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 13;
defparam ram_block1a24.port_b_byte_enable_clock = "clock1";
defparam ram_block1a24.port_b_byte_enable_mask_width = 1;
defparam ram_block1a24.port_b_byte_size = 1;
defparam ram_block1a24.port_b_data_in_clock = "clock1";
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 8191;
defparam ram_block1a24.port_b_logical_ram_depth = 16384;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.port_b_write_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a57(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a57_PORTADATAOUT_bus),
	.portbdataout(ram_block1a57_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena0";
defparam ram_block1a57.clk1_core_clock_enable = "ena1";
defparam ram_block1a57.clk1_input_clock_enable = "ena1";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a57.operation_mode = "bidir_dual_port";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 13;
defparam ram_block1a57.port_a_byte_enable_mask_width = 1;
defparam ram_block1a57.port_a_byte_size = 1;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "none";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 8192;
defparam ram_block1a57.port_a_first_bit_number = 25;
defparam ram_block1a57.port_a_last_address = 16383;
defparam ram_block1a57.port_a_logical_ram_depth = 16384;
defparam ram_block1a57.port_a_logical_ram_width = 32;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.port_b_address_clear = "none";
defparam ram_block1a57.port_b_address_clock = "clock1";
defparam ram_block1a57.port_b_address_width = 13;
defparam ram_block1a57.port_b_byte_enable_clock = "clock1";
defparam ram_block1a57.port_b_byte_enable_mask_width = 1;
defparam ram_block1a57.port_b_byte_size = 1;
defparam ram_block1a57.port_b_data_in_clock = "clock1";
defparam ram_block1a57.port_b_data_out_clear = "none";
defparam ram_block1a57.port_b_data_out_clock = "none";
defparam ram_block1a57.port_b_data_width = 1;
defparam ram_block1a57.port_b_first_address = 8192;
defparam ram_block1a57.port_b_first_bit_number = 25;
defparam ram_block1a57.port_b_last_address = 16383;
defparam ram_block1a57.port_b_logical_ram_depth = 16384;
defparam ram_block1a57.port_b_logical_ram_width = 32;
defparam ram_block1a57.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.port_b_read_enable_clock = "clock1";
defparam ram_block1a57.port_b_write_enable_clock = "clock1";
defparam ram_block1a57.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.clk1_input_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "bidir_dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 16384;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 13;
defparam ram_block1a25.port_b_byte_enable_clock = "clock1";
defparam ram_block1a25.port_b_byte_enable_mask_width = 1;
defparam ram_block1a25.port_b_byte_size = 1;
defparam ram_block1a25.port_b_data_in_clock = "clock1";
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 8191;
defparam ram_block1a25.port_b_logical_ram_depth = 16384;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.port_b_write_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a58(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a58_PORTADATAOUT_bus),
	.portbdataout(ram_block1a58_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena0";
defparam ram_block1a58.clk1_core_clock_enable = "ena1";
defparam ram_block1a58.clk1_input_clock_enable = "ena1";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a58.operation_mode = "bidir_dual_port";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 13;
defparam ram_block1a58.port_a_byte_enable_mask_width = 1;
defparam ram_block1a58.port_a_byte_size = 1;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "none";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 8192;
defparam ram_block1a58.port_a_first_bit_number = 26;
defparam ram_block1a58.port_a_last_address = 16383;
defparam ram_block1a58.port_a_logical_ram_depth = 16384;
defparam ram_block1a58.port_a_logical_ram_width = 32;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.port_b_address_clear = "none";
defparam ram_block1a58.port_b_address_clock = "clock1";
defparam ram_block1a58.port_b_address_width = 13;
defparam ram_block1a58.port_b_byte_enable_clock = "clock1";
defparam ram_block1a58.port_b_byte_enable_mask_width = 1;
defparam ram_block1a58.port_b_byte_size = 1;
defparam ram_block1a58.port_b_data_in_clock = "clock1";
defparam ram_block1a58.port_b_data_out_clear = "none";
defparam ram_block1a58.port_b_data_out_clock = "none";
defparam ram_block1a58.port_b_data_width = 1;
defparam ram_block1a58.port_b_first_address = 8192;
defparam ram_block1a58.port_b_first_bit_number = 26;
defparam ram_block1a58.port_b_last_address = 16383;
defparam ram_block1a58.port_b_logical_ram_depth = 16384;
defparam ram_block1a58.port_b_logical_ram_width = 32;
defparam ram_block1a58.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.port_b_read_enable_clock = "clock1";
defparam ram_block1a58.port_b_write_enable_clock = "clock1";
defparam ram_block1a58.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.clk1_input_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "bidir_dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 16384;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 13;
defparam ram_block1a26.port_b_byte_enable_clock = "clock1";
defparam ram_block1a26.port_b_byte_enable_mask_width = 1;
defparam ram_block1a26.port_b_byte_size = 1;
defparam ram_block1a26.port_b_data_in_clock = "clock1";
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 8191;
defparam ram_block1a26.port_b_logical_ram_depth = 16384;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.port_b_write_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a59(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a59_PORTADATAOUT_bus),
	.portbdataout(ram_block1a59_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena0";
defparam ram_block1a59.clk1_core_clock_enable = "ena1";
defparam ram_block1a59.clk1_input_clock_enable = "ena1";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a59.operation_mode = "bidir_dual_port";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 13;
defparam ram_block1a59.port_a_byte_enable_mask_width = 1;
defparam ram_block1a59.port_a_byte_size = 1;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "none";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 8192;
defparam ram_block1a59.port_a_first_bit_number = 27;
defparam ram_block1a59.port_a_last_address = 16383;
defparam ram_block1a59.port_a_logical_ram_depth = 16384;
defparam ram_block1a59.port_a_logical_ram_width = 32;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.port_b_address_clear = "none";
defparam ram_block1a59.port_b_address_clock = "clock1";
defparam ram_block1a59.port_b_address_width = 13;
defparam ram_block1a59.port_b_byte_enable_clock = "clock1";
defparam ram_block1a59.port_b_byte_enable_mask_width = 1;
defparam ram_block1a59.port_b_byte_size = 1;
defparam ram_block1a59.port_b_data_in_clock = "clock1";
defparam ram_block1a59.port_b_data_out_clear = "none";
defparam ram_block1a59.port_b_data_out_clock = "none";
defparam ram_block1a59.port_b_data_width = 1;
defparam ram_block1a59.port_b_first_address = 8192;
defparam ram_block1a59.port_b_first_bit_number = 27;
defparam ram_block1a59.port_b_last_address = 16383;
defparam ram_block1a59.port_b_logical_ram_depth = 16384;
defparam ram_block1a59.port_b_logical_ram_width = 32;
defparam ram_block1a59.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.port_b_read_enable_clock = "clock1";
defparam ram_block1a59.port_b_write_enable_clock = "clock1";
defparam ram_block1a59.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.clk1_input_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "bidir_dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 16384;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 13;
defparam ram_block1a27.port_b_byte_enable_clock = "clock1";
defparam ram_block1a27.port_b_byte_enable_mask_width = 1;
defparam ram_block1a27.port_b_byte_size = 1;
defparam ram_block1a27.port_b_data_in_clock = "clock1";
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 8191;
defparam ram_block1a27.port_b_logical_ram_depth = 16384;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.port_b_write_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a60(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a60_PORTADATAOUT_bus),
	.portbdataout(ram_block1a60_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena0";
defparam ram_block1a60.clk1_core_clock_enable = "ena1";
defparam ram_block1a60.clk1_input_clock_enable = "ena1";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a60.operation_mode = "bidir_dual_port";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 13;
defparam ram_block1a60.port_a_byte_enable_mask_width = 1;
defparam ram_block1a60.port_a_byte_size = 1;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "none";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 8192;
defparam ram_block1a60.port_a_first_bit_number = 28;
defparam ram_block1a60.port_a_last_address = 16383;
defparam ram_block1a60.port_a_logical_ram_depth = 16384;
defparam ram_block1a60.port_a_logical_ram_width = 32;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.port_b_address_clear = "none";
defparam ram_block1a60.port_b_address_clock = "clock1";
defparam ram_block1a60.port_b_address_width = 13;
defparam ram_block1a60.port_b_byte_enable_clock = "clock1";
defparam ram_block1a60.port_b_byte_enable_mask_width = 1;
defparam ram_block1a60.port_b_byte_size = 1;
defparam ram_block1a60.port_b_data_in_clock = "clock1";
defparam ram_block1a60.port_b_data_out_clear = "none";
defparam ram_block1a60.port_b_data_out_clock = "none";
defparam ram_block1a60.port_b_data_width = 1;
defparam ram_block1a60.port_b_first_address = 8192;
defparam ram_block1a60.port_b_first_bit_number = 28;
defparam ram_block1a60.port_b_last_address = 16383;
defparam ram_block1a60.port_b_logical_ram_depth = 16384;
defparam ram_block1a60.port_b_logical_ram_width = 32;
defparam ram_block1a60.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.port_b_read_enable_clock = "clock1";
defparam ram_block1a60.port_b_write_enable_clock = "clock1";
defparam ram_block1a60.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.clk1_input_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "bidir_dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 16384;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 13;
defparam ram_block1a28.port_b_byte_enable_clock = "clock1";
defparam ram_block1a28.port_b_byte_enable_mask_width = 1;
defparam ram_block1a28.port_b_byte_size = 1;
defparam ram_block1a28.port_b_data_in_clock = "clock1";
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 8191;
defparam ram_block1a28.port_b_logical_ram_depth = 16384;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.port_b_write_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a61(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a61_PORTADATAOUT_bus),
	.portbdataout(ram_block1a61_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena0";
defparam ram_block1a61.clk1_core_clock_enable = "ena1";
defparam ram_block1a61.clk1_input_clock_enable = "ena1";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a61.operation_mode = "bidir_dual_port";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 13;
defparam ram_block1a61.port_a_byte_enable_mask_width = 1;
defparam ram_block1a61.port_a_byte_size = 1;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "none";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 8192;
defparam ram_block1a61.port_a_first_bit_number = 29;
defparam ram_block1a61.port_a_last_address = 16383;
defparam ram_block1a61.port_a_logical_ram_depth = 16384;
defparam ram_block1a61.port_a_logical_ram_width = 32;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.port_b_address_clear = "none";
defparam ram_block1a61.port_b_address_clock = "clock1";
defparam ram_block1a61.port_b_address_width = 13;
defparam ram_block1a61.port_b_byte_enable_clock = "clock1";
defparam ram_block1a61.port_b_byte_enable_mask_width = 1;
defparam ram_block1a61.port_b_byte_size = 1;
defparam ram_block1a61.port_b_data_in_clock = "clock1";
defparam ram_block1a61.port_b_data_out_clear = "none";
defparam ram_block1a61.port_b_data_out_clock = "none";
defparam ram_block1a61.port_b_data_width = 1;
defparam ram_block1a61.port_b_first_address = 8192;
defparam ram_block1a61.port_b_first_bit_number = 29;
defparam ram_block1a61.port_b_last_address = 16383;
defparam ram_block1a61.port_b_logical_ram_depth = 16384;
defparam ram_block1a61.port_b_logical_ram_width = 32;
defparam ram_block1a61.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.port_b_read_enable_clock = "clock1";
defparam ram_block1a61.port_b_write_enable_clock = "clock1";
defparam ram_block1a61.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.clk1_input_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "bidir_dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 16384;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 13;
defparam ram_block1a29.port_b_byte_enable_clock = "clock1";
defparam ram_block1a29.port_b_byte_enable_mask_width = 1;
defparam ram_block1a29.port_b_byte_size = 1;
defparam ram_block1a29.port_b_data_in_clock = "clock1";
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 8191;
defparam ram_block1a29.port_b_logical_ram_depth = 16384;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.port_b_write_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a62(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a62_PORTADATAOUT_bus),
	.portbdataout(ram_block1a62_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena0";
defparam ram_block1a62.clk1_core_clock_enable = "ena1";
defparam ram_block1a62.clk1_input_clock_enable = "ena1";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a62.operation_mode = "bidir_dual_port";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 13;
defparam ram_block1a62.port_a_byte_enable_mask_width = 1;
defparam ram_block1a62.port_a_byte_size = 1;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "none";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 8192;
defparam ram_block1a62.port_a_first_bit_number = 30;
defparam ram_block1a62.port_a_last_address = 16383;
defparam ram_block1a62.port_a_logical_ram_depth = 16384;
defparam ram_block1a62.port_a_logical_ram_width = 32;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.port_b_address_clear = "none";
defparam ram_block1a62.port_b_address_clock = "clock1";
defparam ram_block1a62.port_b_address_width = 13;
defparam ram_block1a62.port_b_byte_enable_clock = "clock1";
defparam ram_block1a62.port_b_byte_enable_mask_width = 1;
defparam ram_block1a62.port_b_byte_size = 1;
defparam ram_block1a62.port_b_data_in_clock = "clock1";
defparam ram_block1a62.port_b_data_out_clear = "none";
defparam ram_block1a62.port_b_data_out_clock = "none";
defparam ram_block1a62.port_b_data_width = 1;
defparam ram_block1a62.port_b_first_address = 8192;
defparam ram_block1a62.port_b_first_bit_number = 30;
defparam ram_block1a62.port_b_last_address = 16383;
defparam ram_block1a62.port_b_logical_ram_depth = 16384;
defparam ram_block1a62.port_b_logical_ram_width = 32;
defparam ram_block1a62.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.port_b_read_enable_clock = "clock1";
defparam ram_block1a62.port_b_write_enable_clock = "clock1";
defparam ram_block1a62.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.clk1_input_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "bidir_dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 16384;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 13;
defparam ram_block1a30.port_b_byte_enable_clock = "clock1";
defparam ram_block1a30.port_b_byte_enable_mask_width = 1;
defparam ram_block1a30.port_b_byte_size = 1;
defparam ram_block1a30.port_b_data_in_clock = "clock1";
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 8191;
defparam ram_block1a30.port_b_logical_ram_depth = 16384;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.port_b_write_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a63(
	.portawe(\decode2|eq_node[1]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a63_PORTADATAOUT_bus),
	.portbdataout(ram_block1a63_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena0";
defparam ram_block1a63.clk1_core_clock_enable = "ena1";
defparam ram_block1a63.clk1_input_clock_enable = "ena1";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a63.operation_mode = "bidir_dual_port";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 13;
defparam ram_block1a63.port_a_byte_enable_mask_width = 1;
defparam ram_block1a63.port_a_byte_size = 1;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "none";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 8192;
defparam ram_block1a63.port_a_first_bit_number = 31;
defparam ram_block1a63.port_a_last_address = 16383;
defparam ram_block1a63.port_a_logical_ram_depth = 16384;
defparam ram_block1a63.port_a_logical_ram_width = 32;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.port_b_address_clear = "none";
defparam ram_block1a63.port_b_address_clock = "clock1";
defparam ram_block1a63.port_b_address_width = 13;
defparam ram_block1a63.port_b_byte_enable_clock = "clock1";
defparam ram_block1a63.port_b_byte_enable_mask_width = 1;
defparam ram_block1a63.port_b_byte_size = 1;
defparam ram_block1a63.port_b_data_in_clock = "clock1";
defparam ram_block1a63.port_b_data_out_clear = "none";
defparam ram_block1a63.port_b_data_out_clock = "none";
defparam ram_block1a63.port_b_data_width = 1;
defparam ram_block1a63.port_b_first_address = 8192;
defparam ram_block1a63.port_b_first_bit_number = 31;
defparam ram_block1a63.port_b_last_address = 16383;
defparam ram_block1a63.port_b_logical_ram_depth = 16384;
defparam ram_block1a63.port_b_logical_ram_width = 32;
defparam ram_block1a63.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.port_b_read_enable_clock = "clock1";
defparam ram_block1a63.port_b_write_enable_clock = "clock1";
defparam ram_block1a63.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(\decode2|eq_node[0]~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.clk1_input_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_m062:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "bidir_dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 16384;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 13;
defparam ram_block1a31.port_b_byte_enable_clock = "clock1";
defparam ram_block1a31.port_b_byte_enable_mask_width = 1;
defparam ram_block1a31.port_b_byte_size = 1;
defparam ram_block1a31.port_b_data_in_clock = "clock1";
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 8191;
defparam ram_block1a31.port_b_logical_ram_depth = 16384;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.port_b_write_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(address_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clocken0),
	.q(address_reg_a_0),
	.prn(vcc));
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";

endmodule

module Computer_System_decode_5la (
	readaddress_15,
	writeaddress_15,
	saved_grant_0,
	saved_grant_1,
	wren,
	eq_node_1,
	eq_node_0)/* synthesis synthesis_greybox=0 */;
input 	readaddress_15;
input 	writeaddress_15;
input 	saved_grant_0;
input 	saved_grant_1;
input 	wren;
output 	eq_node_1;
output 	eq_node_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \eq_node[1] (
	.dataa(!saved_grant_0),
	.datab(!readaddress_15),
	.datac(!saved_grant_1),
	.datad(!writeaddress_15),
	.datae(!wren),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(eq_node_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \eq_node[1] .extended_lut = "off";
defparam \eq_node[1] .lut_mask = 64'h0000111F0000111F;
defparam \eq_node[1] .shared_arith = "off";

cyclonev_lcell_comb \eq_node[0] (
	.dataa(!saved_grant_0),
	.datab(!readaddress_15),
	.datac(!saved_grant_1),
	.datad(!writeaddress_15),
	.datae(!wren),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(eq_node_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \eq_node[0] .extended_lut = "off";
defparam \eq_node[0] .lut_mask = 64'h0000EEE00000EEE0;
defparam \eq_node[0] .shared_arith = "off";

endmodule

module Computer_System_decode_5la_1 (
	eq_node_1,
	eq_node_0,
	onchip_sram_s2_address_13,
	onchip_sram_s2_chipselect,
	onchip_sram_s2_write)/* synthesis synthesis_greybox=0 */;
output 	eq_node_1;
output 	eq_node_0;
input 	onchip_sram_s2_address_13;
input 	onchip_sram_s2_chipselect;
input 	onchip_sram_s2_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \eq_node[1]~0 (
	.dataa(!onchip_sram_s2_address_13),
	.datab(!onchip_sram_s2_chipselect),
	.datac(!onchip_sram_s2_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(eq_node_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \eq_node[1]~0 .extended_lut = "off";
defparam \eq_node[1]~0 .lut_mask = 64'h0101010101010101;
defparam \eq_node[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \eq_node[0]~1 (
	.dataa(!onchip_sram_s2_address_13),
	.datab(!onchip_sram_s2_chipselect),
	.datac(!onchip_sram_s2_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(eq_node_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \eq_node[0]~1 .extended_lut = "off";
defparam \eq_node[0]~1 .lut_mask = 64'h0202020202020202;
defparam \eq_node[0]~1 .shared_arith = "off";

endmodule

module Computer_System_mux_2hb (
	ram_block1a40,
	ram_block1a8,
	ram_block1a41,
	ram_block1a9,
	ram_block1a42,
	ram_block1a10,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a48,
	ram_block1a16,
	ram_block1a49,
	ram_block1a17,
	ram_block1a50,
	ram_block1a18,
	ram_block1a51,
	ram_block1a19,
	ram_block1a52,
	ram_block1a20,
	ram_block1a53,
	ram_block1a21,
	ram_block1a54,
	ram_block1a22,
	ram_block1a55,
	ram_block1a23,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a59,
	ram_block1a27,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	address_reg_a_0,
	l1_w16_n0_mux_dataout,
	l1_w17_n0_mux_dataout,
	l1_w18_n0_mux_dataout,
	l1_w19_n0_mux_dataout,
	l1_w20_n0_mux_dataout,
	l1_w21_n0_mux_dataout,
	l1_w22_n0_mux_dataout,
	l1_w23_n0_mux_dataout,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a40;
input 	ram_block1a8;
input 	ram_block1a41;
input 	ram_block1a9;
input 	ram_block1a42;
input 	ram_block1a10;
input 	ram_block1a43;
input 	ram_block1a11;
input 	ram_block1a44;
input 	ram_block1a12;
input 	ram_block1a45;
input 	ram_block1a13;
input 	ram_block1a46;
input 	ram_block1a14;
input 	ram_block1a47;
input 	ram_block1a15;
input 	ram_block1a48;
input 	ram_block1a16;
input 	ram_block1a49;
input 	ram_block1a17;
input 	ram_block1a50;
input 	ram_block1a18;
input 	ram_block1a51;
input 	ram_block1a19;
input 	ram_block1a52;
input 	ram_block1a20;
input 	ram_block1a53;
input 	ram_block1a21;
input 	ram_block1a54;
input 	ram_block1a22;
input 	ram_block1a55;
input 	ram_block1a23;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	address_reg_a_0;
output 	l1_w16_n0_mux_dataout;
output 	l1_w17_n0_mux_dataout;
output 	l1_w18_n0_mux_dataout;
output 	l1_w19_n0_mux_dataout;
output 	l1_w20_n0_mux_dataout;
output 	l1_w21_n0_mux_dataout;
output 	l1_w22_n0_mux_dataout;
output 	l1_w23_n0_mux_dataout;
output 	l1_w8_n0_mux_dataout;
output 	l1_w9_n0_mux_dataout;
output 	l1_w10_n0_mux_dataout;
output 	l1_w11_n0_mux_dataout;
output 	l1_w12_n0_mux_dataout;
output 	l1_w13_n0_mux_dataout;
output 	l1_w14_n0_mux_dataout;
output 	l1_w15_n0_mux_dataout;
output 	l1_w24_n0_mux_dataout;
output 	l1_w25_n0_mux_dataout;
output 	l1_w26_n0_mux_dataout;
output 	l1_w27_n0_mux_dataout;
output 	l1_w28_n0_mux_dataout;
output 	l1_w29_n0_mux_dataout;
output 	l1_w30_n0_mux_dataout;
output 	l1_w31_n0_mux_dataout;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \l1_w16_n0_mux_dataout~0 (
	.dataa(!ram_block1a48),
	.datab(!ram_block1a16),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w16_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w16_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w16_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w16_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w17_n0_mux_dataout~0 (
	.dataa(!ram_block1a49),
	.datab(!ram_block1a17),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w17_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w17_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w17_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w17_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w18_n0_mux_dataout~0 (
	.dataa(!ram_block1a50),
	.datab(!ram_block1a18),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w18_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w18_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w18_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w18_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w19_n0_mux_dataout~0 (
	.dataa(!ram_block1a51),
	.datab(!ram_block1a19),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w19_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w19_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w19_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w19_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w20_n0_mux_dataout~0 (
	.dataa(!ram_block1a52),
	.datab(!ram_block1a20),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w20_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w20_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w20_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w20_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w21_n0_mux_dataout~0 (
	.dataa(!ram_block1a53),
	.datab(!ram_block1a21),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w21_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w21_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w21_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w21_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w22_n0_mux_dataout~0 (
	.dataa(!ram_block1a54),
	.datab(!ram_block1a22),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w22_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w22_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w22_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w22_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w23_n0_mux_dataout~0 (
	.dataa(!ram_block1a55),
	.datab(!ram_block1a23),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w23_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w23_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w23_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w23_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w8_n0_mux_dataout~0 (
	.dataa(!ram_block1a40),
	.datab(!ram_block1a8),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w8_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w8_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w8_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w8_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w9_n0_mux_dataout~0 (
	.dataa(!ram_block1a41),
	.datab(!ram_block1a9),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w9_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w9_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w9_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w9_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w10_n0_mux_dataout~0 (
	.dataa(!ram_block1a42),
	.datab(!ram_block1a10),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w10_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w10_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w10_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w10_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w11_n0_mux_dataout~0 (
	.dataa(!ram_block1a43),
	.datab(!ram_block1a11),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w11_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w11_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w11_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w11_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w12_n0_mux_dataout~0 (
	.dataa(!ram_block1a44),
	.datab(!ram_block1a12),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w12_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w12_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w12_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w12_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w13_n0_mux_dataout~0 (
	.dataa(!ram_block1a45),
	.datab(!ram_block1a13),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w13_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w13_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w13_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w13_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w14_n0_mux_dataout~0 (
	.dataa(!ram_block1a46),
	.datab(!ram_block1a14),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w14_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w14_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w14_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w14_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w15_n0_mux_dataout~0 (
	.dataa(!ram_block1a47),
	.datab(!ram_block1a15),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w15_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w15_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w15_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w15_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w24_n0_mux_dataout~0 (
	.dataa(!ram_block1a56),
	.datab(!ram_block1a24),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w24_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w24_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w24_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w24_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w25_n0_mux_dataout~0 (
	.dataa(!ram_block1a57),
	.datab(!ram_block1a25),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w25_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w25_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w25_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w25_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w26_n0_mux_dataout~0 (
	.dataa(!ram_block1a58),
	.datab(!ram_block1a26),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w26_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w26_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w26_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w26_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w27_n0_mux_dataout~0 (
	.dataa(!ram_block1a59),
	.datab(!ram_block1a27),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w27_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w27_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w27_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w27_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w28_n0_mux_dataout~0 (
	.dataa(!ram_block1a60),
	.datab(!ram_block1a28),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w28_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w28_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w28_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w28_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w29_n0_mux_dataout~0 (
	.dataa(!ram_block1a61),
	.datab(!ram_block1a29),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w29_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w29_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w29_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w29_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w30_n0_mux_dataout~0 (
	.dataa(!ram_block1a62),
	.datab(!ram_block1a30),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w30_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w30_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w30_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w30_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w31_n0_mux_dataout~0 (
	.dataa(!ram_block1a63),
	.datab(!ram_block1a31),
	.datac(!address_reg_a_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w31_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w31_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w31_n0_mux_dataout~0 .lut_mask = 64'h3535353535353535;
defparam \l1_w31_n0_mux_dataout~0 .shared_arith = "off";

endmodule

module Computer_System_mux_2hb_1 (
	ram_block1a32,
	ram_block1a0,
	ram_block1a33,
	ram_block1a1,
	ram_block1a34,
	ram_block1a2,
	ram_block1a35,
	ram_block1a3,
	ram_block1a36,
	ram_block1a4,
	ram_block1a37,
	ram_block1a5,
	ram_block1a38,
	ram_block1a6,
	ram_block1a39,
	ram_block1a7,
	ram_block1a40,
	ram_block1a8,
	ram_block1a41,
	ram_block1a9,
	ram_block1a42,
	ram_block1a10,
	ram_block1a43,
	ram_block1a11,
	ram_block1a44,
	ram_block1a12,
	ram_block1a45,
	ram_block1a13,
	ram_block1a46,
	ram_block1a14,
	ram_block1a47,
	ram_block1a15,
	ram_block1a48,
	ram_block1a16,
	ram_block1a49,
	ram_block1a17,
	ram_block1a50,
	ram_block1a18,
	ram_block1a51,
	ram_block1a19,
	ram_block1a52,
	ram_block1a20,
	ram_block1a53,
	ram_block1a21,
	ram_block1a54,
	ram_block1a22,
	ram_block1a55,
	ram_block1a23,
	ram_block1a56,
	ram_block1a24,
	ram_block1a57,
	ram_block1a25,
	ram_block1a58,
	ram_block1a26,
	ram_block1a59,
	ram_block1a27,
	ram_block1a60,
	ram_block1a28,
	ram_block1a61,
	ram_block1a29,
	ram_block1a62,
	ram_block1a30,
	ram_block1a63,
	ram_block1a31,
	address_reg_b_0,
	l1_w0_n0_mux_dataout,
	l1_w1_n0_mux_dataout,
	l1_w2_n0_mux_dataout,
	l1_w3_n0_mux_dataout,
	l1_w4_n0_mux_dataout,
	l1_w5_n0_mux_dataout,
	l1_w6_n0_mux_dataout,
	l1_w7_n0_mux_dataout,
	l1_w8_n0_mux_dataout,
	l1_w9_n0_mux_dataout,
	l1_w10_n0_mux_dataout,
	l1_w11_n0_mux_dataout,
	l1_w12_n0_mux_dataout,
	l1_w13_n0_mux_dataout,
	l1_w14_n0_mux_dataout,
	l1_w15_n0_mux_dataout,
	l1_w16_n0_mux_dataout,
	l1_w17_n0_mux_dataout,
	l1_w18_n0_mux_dataout,
	l1_w19_n0_mux_dataout,
	l1_w20_n0_mux_dataout,
	l1_w21_n0_mux_dataout,
	l1_w22_n0_mux_dataout,
	l1_w23_n0_mux_dataout,
	l1_w24_n0_mux_dataout,
	l1_w25_n0_mux_dataout,
	l1_w26_n0_mux_dataout,
	l1_w27_n0_mux_dataout,
	l1_w28_n0_mux_dataout,
	l1_w29_n0_mux_dataout,
	l1_w30_n0_mux_dataout,
	l1_w31_n0_mux_dataout)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a32;
input 	ram_block1a0;
input 	ram_block1a33;
input 	ram_block1a1;
input 	ram_block1a34;
input 	ram_block1a2;
input 	ram_block1a35;
input 	ram_block1a3;
input 	ram_block1a36;
input 	ram_block1a4;
input 	ram_block1a37;
input 	ram_block1a5;
input 	ram_block1a38;
input 	ram_block1a6;
input 	ram_block1a39;
input 	ram_block1a7;
input 	ram_block1a40;
input 	ram_block1a8;
input 	ram_block1a41;
input 	ram_block1a9;
input 	ram_block1a42;
input 	ram_block1a10;
input 	ram_block1a43;
input 	ram_block1a11;
input 	ram_block1a44;
input 	ram_block1a12;
input 	ram_block1a45;
input 	ram_block1a13;
input 	ram_block1a46;
input 	ram_block1a14;
input 	ram_block1a47;
input 	ram_block1a15;
input 	ram_block1a48;
input 	ram_block1a16;
input 	ram_block1a49;
input 	ram_block1a17;
input 	ram_block1a50;
input 	ram_block1a18;
input 	ram_block1a51;
input 	ram_block1a19;
input 	ram_block1a52;
input 	ram_block1a20;
input 	ram_block1a53;
input 	ram_block1a21;
input 	ram_block1a54;
input 	ram_block1a22;
input 	ram_block1a55;
input 	ram_block1a23;
input 	ram_block1a56;
input 	ram_block1a24;
input 	ram_block1a57;
input 	ram_block1a25;
input 	ram_block1a58;
input 	ram_block1a26;
input 	ram_block1a59;
input 	ram_block1a27;
input 	ram_block1a60;
input 	ram_block1a28;
input 	ram_block1a61;
input 	ram_block1a29;
input 	ram_block1a62;
input 	ram_block1a30;
input 	ram_block1a63;
input 	ram_block1a31;
input 	address_reg_b_0;
output 	l1_w0_n0_mux_dataout;
output 	l1_w1_n0_mux_dataout;
output 	l1_w2_n0_mux_dataout;
output 	l1_w3_n0_mux_dataout;
output 	l1_w4_n0_mux_dataout;
output 	l1_w5_n0_mux_dataout;
output 	l1_w6_n0_mux_dataout;
output 	l1_w7_n0_mux_dataout;
output 	l1_w8_n0_mux_dataout;
output 	l1_w9_n0_mux_dataout;
output 	l1_w10_n0_mux_dataout;
output 	l1_w11_n0_mux_dataout;
output 	l1_w12_n0_mux_dataout;
output 	l1_w13_n0_mux_dataout;
output 	l1_w14_n0_mux_dataout;
output 	l1_w15_n0_mux_dataout;
output 	l1_w16_n0_mux_dataout;
output 	l1_w17_n0_mux_dataout;
output 	l1_w18_n0_mux_dataout;
output 	l1_w19_n0_mux_dataout;
output 	l1_w20_n0_mux_dataout;
output 	l1_w21_n0_mux_dataout;
output 	l1_w22_n0_mux_dataout;
output 	l1_w23_n0_mux_dataout;
output 	l1_w24_n0_mux_dataout;
output 	l1_w25_n0_mux_dataout;
output 	l1_w26_n0_mux_dataout;
output 	l1_w27_n0_mux_dataout;
output 	l1_w28_n0_mux_dataout;
output 	l1_w29_n0_mux_dataout;
output 	l1_w30_n0_mux_dataout;
output 	l1_w31_n0_mux_dataout;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \l1_w0_n0_mux_dataout~0 (
	.dataa(!ram_block1a32),
	.datab(!address_reg_b_0),
	.datac(!ram_block1a0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w0_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w0_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w0_n0_mux_dataout~0 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \l1_w0_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w1_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a33),
	.datac(!ram_block1a1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w1_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w1_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w1_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w1_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w2_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a34),
	.datac(!ram_block1a2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w2_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w2_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w2_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w2_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w3_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a35),
	.datac(!ram_block1a3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w3_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w3_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w3_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w3_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w4_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a36),
	.datac(!ram_block1a4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w4_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w4_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w4_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w4_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w5_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a37),
	.datac(!ram_block1a5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w5_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w5_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w5_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w5_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w6_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a38),
	.datac(!ram_block1a6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w6_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w6_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w6_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w6_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w7_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a39),
	.datac(!ram_block1a7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w7_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w7_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w7_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w7_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w8_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a40),
	.datac(!ram_block1a8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w8_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w8_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w8_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w8_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w9_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a41),
	.datac(!ram_block1a9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w9_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w9_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w9_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w9_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w10_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a42),
	.datac(!ram_block1a10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w10_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w10_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w10_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w10_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w11_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a43),
	.datac(!ram_block1a11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w11_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w11_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w11_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w11_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w12_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a44),
	.datac(!ram_block1a12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w12_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w12_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w12_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w12_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w13_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a45),
	.datac(!ram_block1a13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w13_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w13_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w13_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w13_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w14_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a46),
	.datac(!ram_block1a14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w14_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w14_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w14_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w14_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w15_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a47),
	.datac(!ram_block1a15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w15_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w15_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w15_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w15_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w16_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a48),
	.datac(!ram_block1a16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w16_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w16_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w16_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w16_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w17_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a49),
	.datac(!ram_block1a17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w17_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w17_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w17_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w17_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w18_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a50),
	.datac(!ram_block1a18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w18_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w18_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w18_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w18_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w19_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a51),
	.datac(!ram_block1a19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w19_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w19_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w19_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w19_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w20_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a52),
	.datac(!ram_block1a20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w20_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w20_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w20_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w20_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w21_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a53),
	.datac(!ram_block1a21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w21_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w21_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w21_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w21_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w22_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a54),
	.datac(!ram_block1a22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w22_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w22_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w22_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w22_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w23_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a55),
	.datac(!ram_block1a23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w23_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w23_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w23_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w23_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w24_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a56),
	.datac(!ram_block1a24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w24_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w24_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w24_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w24_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w25_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a57),
	.datac(!ram_block1a25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w25_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w25_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w25_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w25_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w26_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a58),
	.datac(!ram_block1a26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w26_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w26_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w26_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w26_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w27_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a59),
	.datac(!ram_block1a27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w27_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w27_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w27_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w27_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w28_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a60),
	.datac(!ram_block1a28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w28_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w28_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w28_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w28_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w29_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a61),
	.datac(!ram_block1a29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w29_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w29_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w29_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w29_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w30_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a62),
	.datac(!ram_block1a30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w30_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w30_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w30_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w30_n0_mux_dataout~0 .shared_arith = "off";

cyclonev_lcell_comb \l1_w31_n0_mux_dataout~0 (
	.dataa(!address_reg_b_0),
	.datab(!ram_block1a63),
	.datac(!ram_block1a31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(l1_w31_n0_mux_dataout),
	.sumout(),
	.cout(),
	.shareout());
defparam \l1_w31_n0_mux_dataout~0 .extended_lut = "off";
defparam \l1_w31_n0_mux_dataout~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \l1_w31_n0_mux_dataout~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_System_PLL (
	outclk_wire_1,
	outclk_wire_0,
	locked_wire_0,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_1;
output 	outclk_wire_0;
output 	locked_wire_0;
input 	system_pll_ref_clk_clk;
input 	system_pll_ref_reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_System_PLL_sys_pll sys_pll(
	.outclk_wire_1(outclk_wire_1),
	.outclk_wire_0(outclk_wire_0),
	.locked(locked_wire_0),
	.system_pll_ref_clk_clk(system_pll_ref_clk_clk),
	.system_pll_ref_reset_reset(system_pll_ref_reset_reset));

endmodule

module Computer_System_Computer_System_System_PLL_sys_pll (
	outclk_wire_1,
	outclk_wire_0,
	locked,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_1;
output 	outclk_wire_0;
output 	locked;
input 	system_pll_ref_clk_clk;
input 	system_pll_ref_reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_pll_1 altera_pll_i(
	.outclk({outclk_wire_1,outclk_wire_0}),
	.locked(locked),
	.refclk(system_pll_ref_clk_clk),
	.rst(system_pll_ref_reset_reset));

endmodule

module Computer_System_altera_pll_1 (
	outclk,
	locked,
	refclk,
	rst)/* synthesis synthesis_greybox=0 */;
output 	[1:0] outclk;
output 	locked;
input 	refclk;
input 	rst;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fboutclk_wire[0] ;


generic_pll \general[1].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[1]),
	.fboutclk(),
	.locked(),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[1].gpll .clock_name_global = "false";
defparam \general[1].gpll .duty_cycle = 50;
defparam \general[1].gpll .fractional_vco_multiplier = "false";
defparam \general[1].gpll .output_clock_frequency = "100.0 mhz";
defparam \general[1].gpll .phase_shift = "-3000 ps";
defparam \general[1].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[1].gpll .simulation_type = "timing";

generic_pll \general[0].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[0]),
	.fboutclk(\fboutclk_wire[0] ),
	.locked(locked),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[0].gpll .clock_name_global = "false";
defparam \general[0].gpll .duty_cycle = 50;
defparam \general[0].gpll .fractional_vco_multiplier = "false";
defparam \general[0].gpll .output_clock_frequency = "100.0 mhz";
defparam \general[0].gpll .phase_shift = "0 ps";
defparam \general[0].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[0].gpll .simulation_type = "timing";

endmodule
